VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__nfet_01v8_648S5X
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__nfet_01v8_648S5X ;
  ORIGIN 0.790 1.285 ;
  SIZE 1.580 BY 2.570 ;
  OBS
      LAYER pwell ;
        RECT -1.055 -1.550 1.055 1.550 ;
      LAYER li1 ;
        RECT -0.875 1.200 0.875 1.370 ;
        RECT -0.875 -1.200 -0.705 1.200 ;
        RECT -0.165 0.690 0.165 0.860 ;
        RECT -0.305 -0.520 -0.135 0.520 ;
        RECT 0.135 -0.520 0.305 0.520 ;
        RECT -0.165 -0.860 0.165 -0.690 ;
        RECT 0.705 -1.200 0.875 1.200 ;
        RECT -0.875 -1.370 0.875 -1.200 ;
      LAYER met1 ;
        RECT -0.145 0.660 0.145 0.890 ;
        RECT -0.335 -0.500 -0.105 0.500 ;
        RECT 0.105 -0.500 0.335 0.500 ;
        RECT -0.145 -0.890 0.145 -0.660 ;
  END
END sky130_fd_pr__nfet_01v8_648S5X
MACRO sky130_fd_pr__pfet_01v8_XJ7KDL
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_XJ7KDL ;
  ORIGIN 0.790 2.080 ;
  SIZE 1.580 BY 4.160 ;
  OBS
      LAYER nwell ;
        RECT -1.055 -2.345 1.055 2.345 ;
      LAYER li1 ;
        RECT -0.875 1.995 0.875 2.165 ;
        RECT -0.875 -1.995 -0.705 1.995 ;
        RECT -0.165 1.485 0.165 1.655 ;
        RECT -0.305 -1.270 -0.135 1.270 ;
        RECT 0.135 -1.270 0.305 1.270 ;
        RECT -0.165 -1.655 0.165 -1.485 ;
        RECT 0.705 -1.995 0.875 1.995 ;
        RECT -0.875 -2.165 0.875 -1.995 ;
      LAYER met1 ;
        RECT -0.145 1.455 0.145 1.685 ;
        RECT -0.335 -1.250 -0.105 1.250 ;
        RECT 0.105 -1.250 0.335 1.250 ;
        RECT -0.145 -1.685 0.145 -1.455 ;
  END
END sky130_fd_pr__pfet_01v8_XJ7KDL
MACRO fd
  CLASS BLOCK ;
  FOREIGN fd ;
  ORIGIN 4.165 4.945 ;
  SIZE 46.585 BY 24.340 ;
  PIN VDD
    ANTENNADIFFAREA 2.676600 ;
    PORT
      LAYER nwell ;
        RECT -1.775 0.680 0.335 5.370 ;
      LAYER li1 ;
        RECT -1.185 5.190 -0.215 5.320 ;
        RECT -1.595 5.020 0.155 5.190 ;
        RECT -1.595 1.030 -1.425 5.020 ;
        RECT -1.025 1.755 -0.855 4.295 ;
        RECT -0.015 1.030 0.155 5.020 ;
        RECT -1.595 0.860 0.155 1.030 ;
      LAYER met1 ;
        RECT -1.265 5.880 -0.265 7.230 ;
        RECT -2.265 5.695 -1.945 5.710 ;
        RECT -1.665 5.695 0.145 5.880 ;
        RECT -2.265 5.465 0.145 5.695 ;
        RECT -2.265 5.450 -1.945 5.465 ;
        RECT -1.665 5.010 0.145 5.465 ;
        RECT -2.265 4.150 -1.945 4.165 ;
        RECT -1.055 4.150 -0.825 4.275 ;
        RECT -2.265 3.920 -0.825 4.150 ;
        RECT -2.265 3.905 -1.945 3.920 ;
        RECT -1.055 1.775 -0.825 3.920 ;
      LAYER met2 ;
        RECT -2.235 5.420 -1.975 5.740 ;
        RECT -2.220 4.195 -1.990 5.420 ;
        RECT -2.235 3.875 -1.975 4.195 ;
    END
    PORT
      LAYER nwell ;
        RECT 2.250 1.110 6.940 3.220 ;
      LAYER li1 ;
        RECT 2.430 2.870 6.760 3.040 ;
        RECT 2.430 1.460 2.600 2.870 ;
        RECT 6.590 2.610 6.760 2.870 ;
        RECT 6.590 1.760 6.825 2.610 ;
        RECT 6.590 1.460 6.760 1.760 ;
        RECT 2.430 1.290 6.760 1.460 ;
      LAYER met1 ;
        RECT 6.545 2.700 7.065 2.870 ;
        RECT 6.545 1.680 7.855 2.700 ;
        RECT 6.545 1.300 7.065 1.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.300 12.900 37.100 13.320 ;
        RECT 36.300 11.900 37.960 12.900 ;
        RECT 36.300 11.620 37.100 11.900 ;
    END
    PORT
      LAYER nwell ;
        RECT 35.560 0.610 37.670 5.300 ;
      LAYER li1 ;
        RECT 36.145 5.120 37.115 5.270 ;
        RECT 35.740 4.950 37.490 5.120 ;
        RECT 35.740 0.960 35.910 4.950 ;
        RECT 36.310 1.685 36.480 4.225 ;
        RECT 37.320 0.960 37.490 4.950 ;
        RECT 35.740 0.790 37.490 0.960 ;
      LAYER met1 ;
        RECT 36.080 5.780 37.080 7.170 ;
        RECT 35.720 5.770 37.560 5.780 ;
        RECT 34.920 5.510 37.560 5.770 ;
        RECT 35.720 4.920 37.560 5.510 ;
        RECT 36.280 3.820 36.510 4.205 ;
        RECT 34.920 3.560 36.510 3.820 ;
        RECT 36.280 1.705 36.510 3.560 ;
      LAYER met2 ;
        RECT 34.950 3.530 35.210 5.800 ;
    END
    PORT
      LAYER nwell ;
        RECT 30.540 0.840 32.650 5.530 ;
      LAYER li1 ;
        RECT 31.140 5.350 32.050 5.510 ;
        RECT 30.720 5.180 32.470 5.350 ;
        RECT 30.720 1.190 30.890 5.180 ;
        RECT 31.140 5.170 32.050 5.180 ;
        RECT 31.290 1.915 31.460 4.455 ;
        RECT 32.300 1.190 32.470 5.180 ;
        RECT 30.720 1.020 32.470 1.190 ;
      LAYER met1 ;
        RECT 30.045 5.800 30.365 5.835 ;
        RECT 31.010 5.830 32.010 7.390 ;
        RECT 30.650 5.800 32.470 5.830 ;
        RECT 30.045 5.610 32.470 5.800 ;
        RECT 30.045 5.575 30.365 5.610 ;
        RECT 30.650 5.140 32.470 5.610 ;
        RECT 30.075 3.685 30.335 3.750 ;
        RECT 31.260 3.685 31.490 4.435 ;
        RECT 30.075 3.495 31.490 3.685 ;
        RECT 30.075 3.430 30.335 3.495 ;
        RECT 31.260 1.935 31.490 3.495 ;
      LAYER met2 ;
        RECT 30.075 5.545 30.335 5.865 ;
        RECT 30.110 3.720 30.300 5.545 ;
        RECT 30.045 3.460 30.365 3.720 ;
    END
    PORT
      LAYER nwell ;
        RECT 21.950 1.590 26.640 3.700 ;
      LAYER li1 ;
        RECT 22.130 3.350 26.460 3.520 ;
        RECT 22.130 1.940 22.300 3.350 ;
        RECT 26.290 3.210 26.460 3.350 ;
        RECT 26.290 2.100 26.570 3.210 ;
        RECT 26.290 1.940 26.460 2.100 ;
        RECT 22.130 1.770 26.460 1.940 ;
      LAYER met1 ;
        RECT 26.290 3.230 27.150 3.510 ;
        RECT 26.290 2.230 27.730 3.230 ;
        RECT 26.290 1.800 27.150 2.230 ;
    END
    PORT
      LAYER nwell ;
        RECT 17.180 0.470 19.290 5.160 ;
      LAYER li1 ;
        RECT 17.690 4.980 18.660 5.120 ;
        RECT 17.360 4.810 19.110 4.980 ;
        RECT 17.360 0.820 17.530 4.810 ;
        RECT 17.930 1.545 18.100 4.085 ;
        RECT 18.940 0.820 19.110 4.810 ;
        RECT 17.360 0.650 19.110 0.820 ;
      LAYER met1 ;
        RECT 17.710 5.690 18.710 6.920 ;
        RECT 17.410 5.490 19.140 5.690 ;
        RECT 17.140 5.230 19.140 5.490 ;
        RECT 17.410 4.830 19.140 5.230 ;
        RECT 17.900 3.800 18.130 4.065 ;
        RECT 16.670 3.780 16.990 3.790 ;
        RECT 17.180 3.780 18.130 3.800 ;
        RECT 16.670 3.560 18.130 3.780 ;
        RECT 16.670 3.540 17.430 3.560 ;
        RECT 16.670 3.530 16.990 3.540 ;
        RECT 17.900 1.565 18.130 3.560 ;
      LAYER met2 ;
        RECT 17.170 5.480 17.430 5.520 ;
        RECT 16.710 5.240 17.430 5.480 ;
        RECT 16.710 3.820 16.950 5.240 ;
        RECT 17.170 5.200 17.430 5.240 ;
        RECT 16.700 3.500 16.960 3.820 ;
    END
    PORT
      LAYER nwell ;
        RECT 11.730 0.480 13.840 5.170 ;
      LAYER li1 ;
        RECT 12.330 4.990 13.270 5.030 ;
        RECT 11.910 4.820 13.660 4.990 ;
        RECT 11.910 0.830 12.080 4.820 ;
        RECT 12.480 1.555 12.650 4.095 ;
        RECT 13.490 0.830 13.660 4.820 ;
        RECT 11.910 0.660 13.660 0.830 ;
      LAYER met1 ;
        RECT 12.310 5.690 13.310 6.730 ;
        RECT 11.460 5.425 11.780 5.450 ;
        RECT 12.030 5.425 13.770 5.690 ;
        RECT 11.460 5.215 13.770 5.425 ;
        RECT 11.460 5.190 11.780 5.215 ;
        RECT 12.030 4.750 13.770 5.215 ;
        RECT 11.460 3.890 11.780 3.915 ;
        RECT 12.450 3.890 12.680 4.075 ;
        RECT 11.460 3.680 12.680 3.890 ;
        RECT 11.460 3.655 11.780 3.680 ;
        RECT 12.450 1.575 12.680 3.680 ;
      LAYER met2 ;
        RECT 11.490 5.160 11.750 5.480 ;
        RECT 11.515 3.945 11.725 5.160 ;
        RECT 11.490 3.625 11.750 3.945 ;
    END
    PORT
      LAYER nwell ;
        RECT 11.560 12.020 16.250 14.130 ;
      LAYER li1 ;
        RECT 11.740 13.780 16.070 13.950 ;
        RECT 11.740 12.370 11.910 13.780 ;
        RECT 15.900 13.460 16.070 13.780 ;
        RECT 15.900 12.710 16.210 13.460 ;
        RECT 15.900 12.370 16.070 12.710 ;
        RECT 11.740 12.200 16.070 12.370 ;
      LAYER met1 ;
        RECT 15.900 13.610 16.490 13.920 ;
        RECT 15.900 12.610 17.380 13.610 ;
        RECT 15.900 12.470 16.490 12.610 ;
    END
  END VDD
  PIN GND
    ANTENNADIFFAREA 1.701000 ;
    PORT
      LAYER pwell ;
        RECT -1.795 -2.950 0.315 0.150 ;
      LAYER li1 ;
        RECT -1.615 -0.200 0.135 -0.030 ;
        RECT -1.615 -2.600 -1.445 -0.200 ;
        RECT -0.605 -1.920 -0.435 -0.880 ;
        RECT -0.035 -2.600 0.135 -0.200 ;
        RECT -1.615 -2.770 0.135 -2.600 ;
        RECT -1.165 -2.830 -0.315 -2.770 ;
      LAYER met1 ;
        RECT -0.635 -1.310 -0.405 -0.900 ;
        RECT -0.635 -1.530 0.355 -1.310 ;
        RECT -0.635 -1.900 -0.405 -1.530 ;
        RECT 0.125 -2.570 0.345 -1.530 ;
        RECT -1.645 -2.890 0.345 -2.570 ;
        RECT -1.645 -3.150 0.135 -2.890 ;
        RECT -1.265 -4.140 -0.265 -3.150 ;
    END
    PORT
      LAYER pwell ;
        RECT 2.990 -1.750 6.090 0.360 ;
      LAYER li1 ;
        RECT 3.170 0.010 5.910 0.180 ;
        RECT 3.170 -0.230 3.340 0.010 ;
        RECT 3.085 -1.090 3.340 -0.230 ;
        RECT 3.170 -1.400 3.340 -1.090 ;
        RECT 5.740 -1.400 5.910 0.010 ;
        RECT 3.170 -1.570 5.910 -1.400 ;
      LAYER met1 ;
        RECT 2.705 -0.100 3.355 0.200 ;
        RECT 1.875 -1.100 3.355 -0.100 ;
        RECT 2.705 -1.570 3.355 -1.100 ;
    END
    PORT
      LAYER pwell ;
        RECT 17.240 -3.120 19.350 -0.020 ;
      LAYER li1 ;
        RECT 17.420 -0.370 19.170 -0.200 ;
        RECT 17.420 -2.770 17.590 -0.370 ;
        RECT 18.430 -2.090 18.600 -1.050 ;
        RECT 19.000 -2.770 19.170 -0.370 ;
        RECT 17.420 -2.940 19.170 -2.770 ;
        RECT 17.745 -3.050 18.835 -2.940 ;
      LAYER met1 ;
        RECT 18.400 -1.440 18.630 -1.070 ;
        RECT 18.400 -1.680 19.310 -1.440 ;
        RECT 18.400 -2.070 18.630 -1.680 ;
        RECT 19.070 -2.770 19.310 -1.680 ;
        RECT 17.335 -3.100 19.310 -2.770 ;
        RECT 17.335 -3.370 19.225 -3.100 ;
        RECT 17.945 -4.190 18.945 -3.370 ;
    END
    PORT
      LAYER pwell ;
        RECT 11.760 -2.740 13.870 0.360 ;
      LAYER li1 ;
        RECT 11.940 0.010 13.690 0.180 ;
        RECT 11.940 -2.390 12.110 0.010 ;
        RECT 12.950 -1.710 13.120 -0.670 ;
        RECT 13.520 -2.390 13.690 0.010 ;
        RECT 11.940 -2.560 13.690 -2.390 ;
        RECT 12.380 -2.630 13.250 -2.560 ;
      LAYER met1 ;
        RECT 12.920 -1.080 13.150 -0.690 ;
        RECT 12.920 -1.280 13.810 -1.080 ;
        RECT 12.920 -1.690 13.150 -1.280 ;
        RECT 13.550 -2.370 13.750 -1.280 ;
        RECT 11.980 -2.570 13.750 -2.370 ;
        RECT 11.980 -3.030 13.740 -2.570 ;
        RECT 12.310 -3.770 13.310 -3.030 ;
    END
    PORT
      LAYER pwell ;
        RECT 32.580 8.430 35.680 10.540 ;
      LAYER li1 ;
        RECT 32.760 10.190 35.500 10.360 ;
        RECT 32.760 9.970 32.930 10.190 ;
        RECT 32.750 9.090 32.950 9.970 ;
        RECT 32.760 8.780 32.930 9.090 ;
        RECT 35.330 8.780 35.500 10.190 ;
        RECT 32.760 8.610 35.500 8.780 ;
      LAYER met1 ;
        RECT 32.610 10.030 33.020 10.370 ;
        RECT 31.680 9.030 33.020 10.030 ;
        RECT 32.610 8.610 33.020 9.030 ;
    END
    PORT
      LAYER pwell ;
        RECT 35.590 -2.780 37.700 0.320 ;
        RECT 35.690 -3.080 37.590 -2.780 ;
      LAYER li1 ;
        RECT 35.770 -0.030 37.520 0.140 ;
        RECT 35.770 -2.430 35.940 -0.030 ;
        RECT 36.780 -1.750 36.950 -0.710 ;
        RECT 37.350 -2.430 37.520 -0.030 ;
        RECT 35.770 -2.600 37.520 -2.430 ;
        RECT 36.205 -2.720 37.065 -2.600 ;
      LAYER met1 ;
        RECT 36.750 -1.460 36.980 -0.730 ;
        RECT 36.750 -1.650 37.650 -1.460 ;
        RECT 36.750 -1.730 36.980 -1.650 ;
        RECT 37.460 -2.450 37.650 -1.650 ;
        RECT 35.690 -2.745 37.650 -2.450 ;
        RECT 35.690 -3.080 37.590 -2.745 ;
        RECT 36.190 -4.260 37.190 -3.080 ;
    END
    PORT
      LAYER pwell ;
        RECT 30.570 -2.480 32.680 0.620 ;
        RECT 30.680 -2.860 32.520 -2.480 ;
      LAYER li1 ;
        RECT 30.750 0.270 32.500 0.440 ;
        RECT 30.750 -2.130 30.920 0.270 ;
        RECT 31.760 -1.450 31.930 -0.410 ;
        RECT 32.330 -2.130 32.500 0.270 ;
        RECT 30.750 -2.300 32.500 -2.130 ;
        RECT 31.205 -2.380 32.035 -2.300 ;
      LAYER met1 ;
        RECT 31.730 -0.860 31.960 -0.430 ;
        RECT 31.690 -1.140 32.800 -0.860 ;
        RECT 31.730 -1.430 31.960 -1.140 ;
        RECT 32.520 -2.080 32.800 -1.140 ;
        RECT 30.680 -2.540 32.800 -2.080 ;
        RECT 30.680 -2.860 32.520 -2.540 ;
        RECT 31.360 -3.660 32.360 -2.860 ;
    END
    PORT
      LAYER pwell ;
        RECT 22.790 -1.170 25.890 0.940 ;
      LAYER li1 ;
        RECT 22.970 0.590 25.710 0.760 ;
        RECT 22.970 0.430 23.140 0.590 ;
        RECT 22.910 -0.540 23.140 0.430 ;
        RECT 22.970 -0.820 23.140 -0.540 ;
        RECT 25.540 -0.820 25.710 0.590 ;
        RECT 22.970 -0.990 25.710 -0.820 ;
      LAYER met1 ;
        RECT 22.580 0.340 23.170 0.790 ;
        RECT 21.840 -0.660 23.170 0.340 ;
        RECT 22.580 -1.010 23.170 -0.660 ;
    END
    PORT
      LAYER pwell ;
        RECT 12.390 9.180 15.490 11.290 ;
      LAYER li1 ;
        RECT 12.570 10.940 15.310 11.110 ;
        RECT 12.570 10.700 12.740 10.940 ;
        RECT 12.370 9.800 12.740 10.700 ;
        RECT 12.570 9.530 12.740 9.800 ;
        RECT 15.140 9.530 15.310 10.940 ;
        RECT 12.570 9.360 15.310 9.530 ;
      LAYER met1 ;
        RECT 12.010 10.790 12.750 11.040 ;
        RECT 11.220 9.790 12.750 10.790 ;
        RECT 12.010 9.450 12.750 9.790 ;
    END
  END GND
  PIN clk
    ANTENNAGATEAREA 0.375000 ;
    PORT
      LAYER li1 ;
        RECT 32.600 12.190 32.770 12.520 ;
        RECT 35.740 12.190 35.910 12.520 ;
      LAYER met1 ;
        RECT 33.770 15.000 34.770 16.030 ;
        RECT 34.060 14.575 34.380 15.000 ;
        RECT 32.475 14.285 35.970 14.575 ;
        RECT 32.475 12.500 32.765 14.285 ;
        RECT 32.475 12.210 32.800 12.500 ;
        RECT 32.475 12.165 32.765 12.210 ;
        RECT 35.650 12.180 35.940 12.860 ;
      LAYER met2 ;
        RECT 35.650 12.745 35.940 14.605 ;
        RECT 35.620 12.455 35.970 12.745 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.940 2.000 3.110 2.330 ;
        RECT 6.080 2.000 6.250 2.330 ;
      LAYER met1 ;
        RECT 4.010 4.670 5.010 5.700 ;
        RECT 4.340 4.050 4.590 4.670 ;
        RECT 6.020 4.050 6.280 4.070 ;
        RECT 2.810 3.750 6.290 4.050 ;
        RECT 2.850 2.310 3.110 3.750 ;
        RECT 2.850 2.020 3.140 2.310 ;
        RECT 2.850 1.960 3.110 2.020 ;
        RECT 6.020 1.980 6.280 3.750 ;
    END
    PORT
      LAYER li1 ;
        RECT 23.480 -0.280 23.650 0.050 ;
        RECT 25.030 -0.280 25.200 0.050 ;
      LAYER met1 ;
        RECT 23.430 -1.300 23.680 0.060 ;
        RECT 25.010 0.030 25.250 0.040 ;
        RECT 25.000 -0.260 25.250 0.030 ;
        RECT 25.000 -0.580 25.260 -0.260 ;
        RECT 25.010 -0.610 25.250 -0.580 ;
        RECT 23.420 -1.560 23.680 -1.300 ;
        RECT 24.970 -1.490 25.290 -1.230 ;
        RECT 23.420 -1.710 23.660 -1.560 ;
        RECT 25.010 -1.710 25.250 -1.490 ;
        RECT 23.420 -1.950 25.250 -1.710 ;
        RECT 23.550 -2.290 25.100 -1.950 ;
        RECT 23.860 -3.170 24.860 -2.290 ;
      LAYER met2 ;
        RECT 24.970 -0.550 25.290 -0.290 ;
        RECT 25.010 -1.200 25.250 -0.550 ;
        RECT 25.000 -1.520 25.260 -1.200 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.080 10.070 13.250 10.400 ;
        RECT 14.630 10.070 14.800 10.400 ;
      LAYER met1 ;
        RECT 13.010 10.380 13.250 10.390 ;
        RECT 13.010 10.090 13.280 10.380 ;
        RECT 13.010 8.990 13.250 10.090 ;
        RECT 14.580 9.930 14.840 10.430 ;
        RECT 14.550 8.990 14.870 9.000 ;
        RECT 13.010 8.750 14.870 8.990 ;
        RECT 13.290 7.420 14.290 8.750 ;
        RECT 14.550 8.740 14.870 8.750 ;
      LAYER met2 ;
        RECT 14.550 9.960 14.870 10.220 ;
        RECT 14.580 8.710 14.840 9.960 ;
    END
    PORT
      LAYER li1 ;
        RECT -0.885 4.510 -0.555 4.680 ;
        RECT -0.885 1.370 -0.555 1.540 ;
        RECT -0.905 -0.710 -0.575 -0.540 ;
        RECT -0.905 -2.260 -0.575 -2.090 ;
      LAYER met1 ;
        RECT -0.865 4.700 -0.575 4.710 ;
        RECT -2.855 4.440 -0.525 4.700 ;
        RECT -4.165 1.340 -3.165 1.810 ;
        RECT -2.855 1.550 -2.595 4.440 ;
        RECT -0.865 1.550 -0.575 1.570 ;
        RECT -2.855 1.340 -0.525 1.550 ;
        RECT -4.165 1.290 -0.525 1.340 ;
        RECT -4.165 1.050 -2.575 1.290 ;
        RECT -4.165 0.780 -3.165 1.050 ;
        RECT -2.855 -0.470 -2.595 1.050 ;
        RECT -2.855 -0.730 -0.515 -0.470 ;
        RECT -2.835 -2.060 -2.575 -0.730 ;
        RECT -0.885 -0.740 -0.595 -0.730 ;
        RECT -2.835 -2.320 -0.575 -2.060 ;
    END
  END clk
  OBS
      LAYER nwell ;
        RECT 31.910 11.300 36.600 13.410 ;
      LAYER li1 ;
        RECT 12.250 12.910 12.420 13.240 ;
        RECT 12.635 13.210 15.175 13.380 ;
        RECT 12.635 12.770 15.175 12.940 ;
        RECT 15.390 12.910 15.560 13.240 ;
        RECT 32.090 13.060 36.420 13.230 ;
        RECT 32.090 11.650 32.260 13.060 ;
        RECT 32.985 12.490 35.525 12.660 ;
        RECT 32.985 12.050 35.525 12.220 ;
        RECT 36.250 11.650 36.420 13.060 ;
        RECT 32.090 11.480 36.420 11.650 ;
        RECT 13.420 10.370 14.460 10.540 ;
        RECT 13.420 9.930 14.460 10.100 ;
        RECT 33.270 9.320 33.440 9.650 ;
        RECT 33.610 9.620 34.650 9.790 ;
        RECT 33.610 9.180 34.650 9.350 ;
        RECT 34.820 9.320 34.990 9.650 ;
        RECT 31.430 4.670 31.760 4.840 ;
        RECT 12.620 4.310 12.950 4.480 ;
        RECT 18.070 4.300 18.400 4.470 ;
        RECT -0.585 1.755 -0.415 4.295 ;
        RECT 3.325 2.300 5.865 2.470 ;
        RECT 3.325 1.860 5.865 2.030 ;
        RECT 12.920 1.555 13.090 4.095 ;
        RECT 18.370 1.545 18.540 4.085 ;
        RECT 22.640 2.480 22.810 2.810 ;
        RECT 23.025 2.780 25.565 2.950 ;
        RECT 23.025 2.340 25.565 2.510 ;
        RECT 25.780 2.480 25.950 2.810 ;
        RECT 31.730 1.915 31.900 4.455 ;
        RECT 36.450 4.440 36.780 4.610 ;
        RECT 31.430 1.530 31.760 1.700 ;
        RECT 36.750 1.685 36.920 4.225 ;
        RECT 12.620 1.170 12.950 1.340 ;
        RECT 18.070 1.160 18.400 1.330 ;
        RECT 36.450 1.300 36.780 1.470 ;
        RECT 23.820 0.020 24.860 0.190 ;
        RECT 31.460 -0.240 31.790 -0.070 ;
        RECT 3.680 -0.860 3.850 -0.530 ;
        RECT 4.020 -0.560 5.060 -0.390 ;
        RECT 12.650 -0.500 12.980 -0.330 ;
        RECT 23.820 -0.420 24.860 -0.250 ;
        RECT -1.045 -1.920 -0.875 -0.880 ;
        RECT 4.020 -1.000 5.060 -0.830 ;
        RECT 5.230 -0.860 5.400 -0.530 ;
        RECT 12.510 -1.710 12.680 -0.670 ;
        RECT 18.130 -0.880 18.460 -0.710 ;
        RECT 12.650 -2.050 12.980 -1.880 ;
        RECT 17.990 -2.090 18.160 -1.050 ;
        RECT 31.320 -1.450 31.490 -0.410 ;
        RECT 36.480 -0.540 36.810 -0.370 ;
        RECT 31.460 -1.790 31.790 -1.620 ;
        RECT 36.340 -1.750 36.510 -0.710 ;
        RECT 36.480 -2.090 36.810 -1.920 ;
        RECT 18.130 -2.430 18.460 -2.260 ;
      LAYER met1 ;
        RECT 10.680 19.325 14.180 19.395 ;
        RECT 10.680 19.125 40.750 19.325 ;
        RECT 10.680 12.595 10.950 19.125 ;
        RECT 13.805 19.055 40.750 19.125 ;
        RECT 13.670 15.050 13.980 15.480 ;
        RECT 15.345 15.050 15.605 15.110 ;
        RECT 12.220 14.850 15.605 15.050 ;
        RECT 12.220 13.220 12.420 14.850 ;
        RECT 13.670 14.840 13.980 14.850 ;
        RECT 15.345 14.790 15.605 14.850 ;
        RECT 14.430 14.300 17.750 14.500 ;
        RECT 14.430 13.410 14.630 14.300 ;
        RECT 12.220 12.930 12.450 13.220 ;
        RECT 12.655 13.180 15.155 13.410 ;
        RECT 15.345 13.310 15.605 13.610 ;
        RECT 12.220 12.920 12.420 12.930 ;
        RECT 12.655 12.740 15.155 12.970 ;
        RECT 15.310 12.880 15.640 13.310 ;
        RECT 17.550 13.190 17.750 14.300 ;
        RECT 34.900 13.530 38.500 13.750 ;
        RECT 17.535 12.930 20.465 13.190 ;
        RECT 1.630 12.325 10.950 12.595 ;
        RECT -0.615 3.020 -0.385 4.275 ;
        RECT -0.615 2.810 0.895 3.020 ;
        RECT -0.615 1.775 -0.385 2.810 ;
        RECT 0.640 0.920 0.850 2.810 ;
        RECT 0.635 0.630 1.420 0.920 ;
        RECT 1.630 0.665 1.900 12.325 ;
        RECT 13.750 11.640 13.930 12.740 ;
        RECT 17.550 11.880 17.750 12.930 ;
        RECT 15.800 11.870 17.750 11.880 ;
        RECT 9.695 11.460 13.930 11.640 ;
        RECT 15.590 11.680 17.750 11.870 ;
        RECT 15.590 11.530 15.860 11.680 ;
        RECT 6.630 3.500 6.890 3.560 ;
        RECT 6.630 3.300 8.470 3.500 ;
        RECT 6.630 3.240 6.890 3.300 ;
        RECT 5.280 2.650 5.540 2.970 ;
        RECT 5.310 2.500 5.510 2.650 ;
        RECT 3.345 2.270 5.845 2.500 ;
        RECT 3.345 1.830 5.845 2.060 ;
        RECT 4.420 0.675 4.610 1.830 ;
        RECT 2.165 0.665 4.615 0.675 ;
        RECT -1.835 0.415 -1.515 0.440 ;
        RECT 0.640 0.415 0.850 0.630 ;
        RECT -1.835 0.205 0.850 0.415 ;
        RECT 1.630 0.410 4.615 0.665 ;
        RECT 8.270 0.640 8.470 3.300 ;
        RECT 9.695 0.640 9.875 11.460 ;
        RECT 13.750 10.570 13.930 11.460 ;
        RECT 13.440 10.340 14.440 10.570 ;
        RECT 13.440 9.900 14.440 10.130 ;
        RECT 13.850 9.710 14.050 9.900 ;
        RECT 15.610 9.710 15.810 11.530 ;
        RECT 13.850 9.510 15.810 9.710 ;
        RECT 12.640 4.490 12.930 4.510 ;
        RECT 10.960 4.250 12.930 4.490 ;
        RECT 16.205 4.270 18.465 4.570 ;
        RECT 10.960 1.380 11.240 4.250 ;
        RECT 12.890 2.690 13.120 4.075 ;
        RECT 12.890 2.530 14.120 2.690 ;
        RECT 12.890 1.575 13.120 2.530 ;
        RECT 10.960 1.140 12.980 1.380 ;
        RECT 10.960 0.640 11.240 1.140 ;
        RECT 13.960 0.820 14.120 2.530 ;
        RECT 16.205 1.390 16.505 4.270 ;
        RECT 18.340 2.570 18.570 4.065 ;
        RECT 18.340 2.360 19.785 2.570 ;
        RECT 18.340 1.565 18.570 2.360 ;
        RECT 16.205 1.090 18.425 1.390 ;
        RECT 16.205 0.910 16.505 1.090 ;
        RECT 16.085 0.880 16.505 0.910 ;
        RECT 14.785 0.820 16.505 0.880 ;
        RECT 1.630 0.395 2.340 0.410 ;
        RECT -1.835 0.180 -1.515 0.205 ;
        RECT 4.420 -0.360 4.610 0.410 ;
        RECT 8.255 0.400 11.240 0.640 ;
        RECT 13.950 0.630 16.505 0.820 ;
        RECT 13.950 0.580 15.300 0.630 ;
        RECT 6.480 0.200 8.470 0.400 ;
        RECT 9.695 0.390 9.875 0.400 ;
        RECT 3.645 -0.550 3.835 -0.525 ;
        RECT 3.645 -0.840 3.880 -0.550 ;
        RECT 4.040 -0.590 5.040 -0.360 ;
        RECT -1.835 -1.315 -1.515 -1.290 ;
        RECT -1.075 -1.315 -0.845 -0.900 ;
        RECT -1.835 -1.525 -0.845 -1.315 ;
        RECT -1.835 -1.550 -1.515 -1.525 ;
        RECT -1.075 -1.900 -0.845 -1.525 ;
        RECT 3.645 -1.995 3.835 -0.840 ;
        RECT 4.040 -1.030 5.040 -0.800 ;
        RECT 5.200 -0.820 5.430 -0.550 ;
        RECT 4.470 -1.400 4.670 -1.030 ;
        RECT 5.185 -1.140 5.445 -0.820 ;
        RECT 6.480 -1.060 6.680 0.200 ;
        RECT 10.960 -0.240 11.240 0.400 ;
        RECT 11.920 0.430 12.240 0.480 ;
        RECT 13.960 0.430 14.120 0.580 ;
        RECT 11.920 0.270 14.120 0.430 ;
        RECT 14.785 0.400 15.300 0.580 ;
        RECT 11.920 0.220 12.240 0.270 ;
        RECT 10.960 -0.480 12.990 -0.240 ;
        RECT 10.980 -0.520 12.990 -0.480 ;
        RECT 6.480 -1.150 6.690 -1.060 ;
        RECT 6.490 -1.400 6.690 -1.150 ;
        RECT 4.470 -1.600 6.690 -1.400 ;
        RECT 10.990 -1.840 11.280 -0.520 ;
        RECT 12.670 -0.530 12.960 -0.520 ;
        RECT 11.920 -1.030 12.240 -0.980 ;
        RECT 12.480 -1.030 12.710 -0.690 ;
        RECT 11.920 -1.190 12.710 -1.030 ;
        RECT 11.920 -1.240 12.240 -1.190 ;
        RECT 12.480 -1.690 12.710 -1.190 ;
        RECT 5.185 -1.995 5.445 -1.930 ;
        RECT 3.645 -2.185 5.445 -1.995 ;
        RECT 10.990 -2.120 13.010 -1.840 ;
        RECT 4.440 -2.810 4.660 -2.185 ;
        RECT 5.185 -2.250 5.445 -2.185 ;
        RECT 15.050 -4.695 15.300 0.400 ;
        RECT 16.205 -0.620 16.505 0.630 ;
        RECT 19.570 0.670 19.780 2.360 ;
        RECT 20.205 0.670 20.465 12.930 ;
        RECT 34.900 12.690 35.120 13.530 ;
        RECT 38.280 12.705 38.500 13.530 ;
        RECT 33.005 12.460 35.505 12.690 ;
        RECT 38.280 12.435 40.050 12.705 ;
        RECT 33.005 12.020 35.505 12.250 ;
        RECT 34.040 11.050 34.240 12.020 ;
        RECT 28.885 10.850 34.240 11.050 ;
        RECT 38.280 11.000 38.500 12.435 ;
        RECT 24.000 4.630 24.310 5.270 ;
        RECT 22.600 4.330 26.050 4.630 ;
        RECT 22.600 2.470 22.900 4.330 ;
        RECT 25.300 3.820 28.070 4.000 ;
        RECT 25.300 2.980 25.480 3.820 ;
        RECT 23.045 2.750 25.545 2.980 ;
        RECT 23.045 2.310 25.545 2.540 ;
        RECT 25.720 2.500 26.020 3.060 ;
        RECT 23.950 1.215 24.130 2.310 ;
        RECT 27.890 1.630 28.070 3.820 ;
        RECT 28.885 1.630 29.085 10.850 ;
        RECT 34.040 9.820 34.240 10.850 ;
        RECT 35.890 10.780 38.500 11.000 ;
        RECT 33.260 9.630 33.465 9.680 ;
        RECT 33.240 9.340 33.470 9.630 ;
        RECT 33.630 9.590 34.630 9.820 ;
        RECT 33.260 8.320 33.465 9.340 ;
        RECT 33.630 9.150 34.630 9.380 ;
        RECT 34.080 8.870 34.300 9.150 ;
        RECT 34.780 9.040 35.060 9.650 ;
        RECT 35.890 8.870 36.110 10.780 ;
        RECT 34.080 8.650 36.110 8.870 ;
        RECT 33.220 8.040 35.090 8.320 ;
        RECT 33.900 7.400 34.250 8.040 ;
        RECT 29.665 4.590 31.745 4.870 ;
        RECT 29.665 3.920 29.945 4.590 ;
        RECT 34.300 4.480 36.820 4.780 ;
        RECT 29.665 3.290 29.905 3.920 ;
        RECT 29.665 1.710 29.945 3.290 ;
        RECT 31.700 3.230 31.930 4.435 ;
        RECT 34.300 3.340 34.600 4.480 ;
        RECT 36.470 4.410 36.760 4.480 ;
        RECT 31.700 2.980 33.010 3.230 ;
        RECT 34.300 3.040 35.330 3.340 ;
        RECT 31.700 1.935 31.930 2.980 ;
        RECT 31.450 1.710 31.740 1.730 ;
        RECT 29.665 1.630 31.815 1.710 ;
        RECT 27.880 1.450 31.815 1.630 ;
        RECT 26.110 1.430 31.815 1.450 ;
        RECT 26.110 1.400 30.015 1.430 ;
        RECT 26.110 1.270 28.070 1.400 ;
        RECT 19.570 0.410 20.465 0.670 ;
        RECT 21.310 0.965 24.160 1.215 ;
        RECT 17.385 0.285 17.705 0.310 ;
        RECT 19.570 0.285 19.780 0.410 ;
        RECT 17.385 0.075 19.780 0.285 ;
        RECT 17.385 0.050 17.705 0.075 ;
        RECT 16.205 -0.920 18.525 -0.620 ;
        RECT 16.205 -2.230 16.505 -0.920 ;
        RECT 17.385 -1.395 17.705 -1.370 ;
        RECT 17.960 -1.395 18.190 -1.070 ;
        RECT 17.385 -1.605 18.190 -1.395 ;
        RECT 17.385 -1.630 17.705 -1.605 ;
        RECT 17.960 -2.070 18.190 -1.605 ;
        RECT 16.205 -2.530 18.515 -2.230 ;
        RECT 21.310 -4.695 21.560 0.965 ;
        RECT 23.950 0.220 24.130 0.965 ;
        RECT 23.840 -0.010 24.840 0.220 ;
        RECT 23.840 -0.450 24.840 -0.220 ;
        RECT 24.230 -0.850 24.410 -0.450 ;
        RECT 26.110 -0.850 26.290 1.270 ;
        RECT 24.230 -1.030 26.290 -0.850 ;
        RECT 29.665 0.050 29.945 1.400 ;
        RECT 32.755 1.350 33.005 2.980 ;
        RECT 35.030 1.530 35.330 3.040 ;
        RECT 36.720 2.940 36.950 4.205 ;
        RECT 36.720 2.680 38.220 2.940 ;
        RECT 36.720 1.705 36.950 2.680 ;
        RECT 35.020 1.420 36.840 1.530 ;
        RECT 34.280 1.350 36.840 1.420 ;
        RECT 32.755 1.230 36.840 1.350 ;
        RECT 32.755 1.150 35.330 1.230 ;
        RECT 32.755 1.120 34.530 1.150 ;
        RECT 30.450 0.865 30.770 0.870 ;
        RECT 32.755 0.865 33.005 1.120 ;
        RECT 30.450 0.615 33.005 0.865 ;
        RECT 30.450 0.610 30.770 0.615 ;
        RECT 29.665 -0.230 31.795 0.050 ;
        RECT 29.665 -1.610 29.945 -0.230 ;
        RECT 31.480 -0.270 31.770 -0.230 ;
        RECT 30.480 -0.825 30.740 -0.790 ;
        RECT 31.290 -0.825 31.520 -0.430 ;
        RECT 30.480 -1.075 31.520 -0.825 ;
        RECT 30.480 -1.110 30.740 -1.075 ;
        RECT 31.290 -1.430 31.520 -1.075 ;
        RECT 31.480 -1.610 31.770 -1.590 ;
        RECT 29.665 -1.820 31.770 -1.610 ;
        RECT 29.665 -1.890 31.755 -1.820 ;
        RECT 15.050 -4.945 21.560 -4.695 ;
        RECT 33.765 -4.520 33.985 1.120 ;
        RECT 35.020 -0.270 35.320 1.150 ;
        RECT 37.960 1.110 38.220 2.680 ;
        RECT 39.780 1.110 40.050 12.435 ;
        RECT 40.480 1.110 40.750 19.055 ;
        RECT 37.960 0.840 42.420 1.110 ;
        RECT 37.960 0.630 38.220 0.840 ;
        RECT 35.590 0.370 38.220 0.630 ;
        RECT 39.195 -0.250 41.605 -0.030 ;
        RECT 34.950 -0.340 36.780 -0.270 ;
        RECT 34.950 -0.570 36.790 -0.340 ;
        RECT 35.020 -1.890 35.320 -0.570 ;
        RECT 36.310 -1.110 36.540 -0.730 ;
        RECT 35.590 -1.370 36.540 -1.110 ;
        RECT 36.310 -1.730 36.540 -1.370 ;
        RECT 35.020 -1.900 36.100 -1.890 ;
        RECT 36.500 -1.900 36.790 -1.890 ;
        RECT 35.020 -2.140 36.850 -1.900 ;
        RECT 39.195 -4.520 39.415 -0.250 ;
        RECT 33.765 -4.740 39.415 -4.520 ;
      LAYER met2 ;
        RECT 15.315 14.820 15.635 15.080 ;
        RECT 15.375 13.580 15.575 14.820 ;
        RECT 15.315 13.320 15.635 13.580 ;
        RECT 34.750 9.070 35.090 9.350 ;
        RECT 34.780 8.010 35.060 9.070 ;
        RECT 6.600 3.500 6.920 3.530 ;
        RECT 5.310 3.300 6.920 3.500 ;
        RECT 5.310 2.940 5.510 3.300 ;
        RECT 6.600 3.270 6.920 3.300 ;
        RECT 25.720 3.030 26.020 4.660 ;
        RECT 5.250 2.680 5.570 2.940 ;
        RECT 25.690 2.730 26.050 3.030 ;
        RECT 30.480 0.580 30.740 0.900 ;
        RECT -1.805 0.150 -1.545 0.470 ;
        RECT 11.950 0.190 12.210 0.510 ;
        RECT -1.780 -1.260 -1.570 0.150 ;
        RECT 5.155 -1.110 5.475 -0.850 ;
        RECT 12.000 -0.950 12.160 0.190 ;
        RECT 17.415 0.020 17.675 0.340 ;
        RECT -1.805 -1.580 -1.545 -1.260 ;
        RECT 5.220 -1.960 5.410 -1.110 ;
        RECT 11.950 -1.270 12.210 -0.950 ;
        RECT 17.440 -1.340 17.650 0.020 ;
        RECT 30.485 -0.820 30.735 0.580 ;
        RECT 30.450 -1.080 30.770 -0.820 ;
        RECT 17.415 -1.660 17.675 -1.340 ;
        RECT 35.620 -1.400 35.880 0.660 ;
        RECT 5.155 -2.220 5.475 -1.960 ;
  END
END fd
END LIBRARY

