magic
tech sky130A
magscale 1 2
timestamp 1714651723
<< metal1 >>
rect 3510 10222 13333 10276
rect 3510 7764 3564 10222
rect 13279 9185 13333 10222
rect 13279 9119 13477 9185
rect 13543 9119 13549 9185
rect 3418 7564 3618 7764
rect 3502 7392 3562 7564
rect 13279 7333 13333 9119
rect 2280 6202 2480 6402
rect 2752 6294 2912 6342
rect 2344 6056 2384 6202
rect 12588 6182 12764 6226
rect 12588 6034 12632 6182
rect 11926 5990 12632 6034
rect 21724 5916 21922 5960
rect 21878 5748 21922 5916
rect 3488 5146 3544 5314
rect 3412 4946 3612 5146
rect 3478 4786 3542 4946
rect 13284 4786 13348 5252
rect 3478 4722 16884 4786
rect 16820 4088 16884 4722
rect 8252 3370 8452 3570
rect 21876 3214 21928 5748
rect 17404 3162 21928 3214
rect 17875 2931 17941 2937
rect 16782 1801 16848 2082
rect 17875 1801 17941 2865
rect 16782 1735 17941 1801
rect 16782 1728 16848 1735
<< via1 >>
rect 13477 9119 13543 9185
rect 17875 2865 17941 2931
<< metal2 >>
rect 13477 9185 13543 9191
rect 13543 9119 17941 9185
rect 13477 9113 13543 9119
rect 17875 2931 17941 9119
rect 17869 2865 17875 2931
rect 17941 2865 17947 2931
use fd  x1
timestamp 1713507270
transform -1 0 16679 0 -1 3417
box -833 -989 8484 3879
use fd  x2
timestamp 1713507270
transform 1 0 13456 0 1 5966
box -833 -989 8484 3879
use fd  x3
timestamp 1713507270
transform 1 0 3669 0 1 6040
box -833 -989 8484 3879
<< labels >>
flabel metal1 8252 3370 8452 3570 0 FreeSans 256 0 0 0 f_out
port 2 nsew
flabel metal1 2772 6320 2772 6320 0 FreeSans 256 180 0 0 k
flabel metal1 2366 6090 2366 6090 0 FreeSans 256 0 0 0 k
flabel metal1 2280 6202 2480 6402 0 FreeSans 256 0 0 0 clk1
port 1 nsew
flabel metal1 3412 4946 3612 5146 0 FreeSans 256 0 0 0 GND
port 3 nsew
flabel metal1 3418 7564 3618 7764 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
