* NGSPICE file created from pll.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt pfd_lay f_clk_in VPWR f_vco x13/Y sky130_fd_sc_hd__inv_1_3/Y VGND
Xx1 x9/A x5/C test2 x6/Y VGND VGND VPWR VPWR x9/B sky130_fd_sc_hd__nand4_1
Xx3 f_vco VGND VGND VPWR VPWR x6/B sky130_fd_sc_hd__inv_1
Xx2 x9/B x5/C VGND VGND VPWR VPWR x2/Y sky130_fd_sc_hd__nand2_1
Xx5 x9/B x5/B x5/C VGND VGND VPWR VPWR x6/A sky130_fd_sc_hd__nand3_1
Xx6 x6/A x6/B VGND VGND VPWR VPWR x6/Y sky130_fd_sc_hd__nand2_1
Xx8 test2 x9/Y VGND VGND VPWR VPWR x9/A sky130_fd_sc_hd__nand2_1
Xx9 x9/A x9/B VGND VGND VPWR VPWR x9/Y sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand3_1_0 x9/B test4 x9/A VGND VGND VPWR VPWR sky130_fd_sc_hd__inv_1_3/A
+ sky130_fd_sc_hd__nand3_1
Xx10 x6/Y VGND VGND VPWR VPWR x12/A sky130_fd_sc_hd__inv_1
Xx11 x2/Y x6/Y VGND VGND VPWR VPWR x5/C sky130_fd_sc_hd__nand2_1
Xx12 x12/A VGND VGND VPWR VPWR x5/B sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__inv_1_3/A test1 VGND VGND VPWR VPWR test2
+ sky130_fd_sc_hd__nand2_1
Xx13 x6/A VGND VGND VPWR VPWR x13/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_1/Y VGND VGND VPWR VPWR test4 sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 test2 VGND VGND VPWR VPWR sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_2 f_clk_in VGND VGND VPWR VPWR test1 sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__inv_1_3/Y
+ sky130_fd_sc_hd__inv_1
.ends

.subckt sky130_fd_pr__pfet_01v8_KZR7FM a_18_n54# w_n214_n273# a_n76_n54# a_n33_n151#
X0 a_18_n54# a_n33_n151# a_n76_n54# w_n214_n273# sky130_fd_pr__pfet_01v8 ad=0.1566 pd=1.66 as=0.1566 ps=1.66 w=0.54 l=0.18
.ends

.subckt sky130_fd_pr__pfet_01v8_K9S7EM a_18_n54# w_n214_n273# a_n76_n54# a_n33_n151#
X0 a_18_n54# a_n33_n151# a_n76_n54# w_n214_n273# sky130_fd_pr__pfet_01v8 ad=0.1566 pd=1.66 as=0.1566 ps=1.66 w=0.54 l=0.18
.ends

.subckt sky130_fd_pr__nfet_01v8_6FB46G a_18_n42# a_n33_n130# a_n76_n42# a_n178_n216#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n178_n216# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.18
.ends

.subckt sky130_fd_pr__res_generic_po_447X6E a_n48_165# a_n48_n595#
R0 a_n48_165# a_n48_n595# sky130_fd_pr__res_generic_po w=0.48 l=1.65
.ends

.subckt sky130_fd_pr__pfet_01v8_XJ7KDL w_n211_n469# a_n73_n250# a_n33_n347# a_15_n250#
X0 a_15_n250# a_n33_n347# a_n73_n250# w_n211_n469# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt fd VDD GND clk m1_6090_122#
XXM12 VDD VDD m1_2384_n248# m1_2770_1902# sky130_fd_pr__pfet_01v8_XJ7KDL
XXM14 VDD VDD m1_6090_122# q_b sky130_fd_pr__pfet_01v8_XJ7KDL
XXM13 m1_6090_122# m1_4846_n206# GND GND sky130_fd_pr__nfet_01v8_648S5X
XXM15 m1_2770_1902# m1_2384_n248# GND GND sky130_fd_pr__nfet_01v8_648S5X
XXM16 VDD VDD clk clk_b sky130_fd_pr__pfet_01v8_XJ7KDL
XXM17 VDD VDD m1_4846_n206# m1_6090_122# sky130_fd_pr__pfet_01v8_XJ7KDL
XXM18 clk_b clk GND GND sky130_fd_pr__nfet_01v8_648S5X
XXM1 VDD VDD m1_992_n194# m1_2384_n248# sky130_fd_pr__pfet_01v8_XJ7KDL
XXM2 q_b m1_6090_122# GND GND sky130_fd_pr__nfet_01v8_648S5X
XXM3 XM3/w_n211_n469# m1_4846_n206# clk q_b sky130_fd_pr__pfet_01v8_XJ7KDL
XXM4 m1_4846_n206# clk m1_2384_n248# GND sky130_fd_pr__nfet_01v8_648S5X
XXM5 m1_2384_n248# m1_992_n194# GND GND sky130_fd_pr__nfet_01v8_648S5X
XXM6 VDD q_b clk m1_992_n194# sky130_fd_pr__pfet_01v8_XJ7KDL
XXM7 VDD m1_2770_1902# clk_b m1_992_n194# sky130_fd_pr__pfet_01v8_XJ7KDL
XXM8 m1_2770_1902# clk m1_992_n194# GND sky130_fd_pr__nfet_01v8_648S5X
XXM9 VDD m1_4846_n206# clk_b m1_2384_n248# sky130_fd_pr__pfet_01v8_XJ7KDL
XXM10 q_b clk_b m1_4846_n206# GND sky130_fd_pr__nfet_01v8_648S5X
XXM11 m1_992_n194# clk_b q_b GND sky130_fd_pr__nfet_01v8_648S5X
.ends

.subckt fd_8 VDD k f_out GND
Xx1 VDD GND x1/clk f_out fd
Xx2 VDD GND x2/clk x1/clk fd
Xx3 VDD GND k x2/clk fd
.ends

.subckt sky130_fd_pr__nfet_01v8_HAAXKC a_n76_n1500# a_n33_n1588# a_18_n1500# a_n178_n1674#
X0 a_18_n1500# a_n33_n1588# a_n76_n1500# a_n178_n1674# sky130_fd_pr__nfet_01v8 ad=4.35 pd=30.58 as=4.35 ps=30.58 w=15 l=0.18
.ends

.subckt sky130_fd_pr__pfet_01v8_7PMXFU a_n76_n4500# w_n214_n4719# a_18_n4500# a_n33_n4597#
X0 a_18_n4500# a_n33_n4597# a_n76_n4500# w_n214_n4719# sky130_fd_pr__pfet_01v8 ad=13.05 pd=90.58 as=13.05 ps=90.58 w=45 l=0.18
.ends

.subckt sky130_fd_pr__nfet_01v8_6FB27G a_18_n42# a_n33_n130# a_n76_n42# a_n178_n216#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n178_n216# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.18
.ends

.subckt sky130_fd_pr__pfet_01v8_KXJ7FM a_18_n54# w_n214_n273# a_n76_n54# a_n33_n151#
X0 a_18_n54# a_n33_n151# a_n76_n54# w_n214_n273# sky130_fd_pr__pfet_01v8 ad=0.1566 pd=1.66 as=0.1566 ps=1.66 w=0.54 l=0.18
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_39XMLG m3_10038_n15680# c1_n3146_n15640# c1_10078_n15640#
+ c1_3466_n15640# c1_n16370_n15640# m3_n9798_n15680# m3_n3186_n15680# c1_n9758_n15640#
+ m3_3426_n15680# m3_n16410_n15680#
X0 c1_n16370_n15640# m3_n16410_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X1 c1_n3146_n15640# m3_n3186_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X2 c1_n3146_n15640# m3_n3186_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X3 c1_3466_n15640# m3_3426_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X4 c1_3466_n15640# m3_3426_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X5 c1_3466_n15640# m3_3426_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X6 c1_n16370_n15640# m3_n16410_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X7 c1_n16370_n15640# m3_n16410_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X8 c1_3466_n15640# m3_3426_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X9 c1_n3146_n15640# m3_n3186_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X10 c1_10078_n15640# m3_10038_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X11 c1_10078_n15640# m3_10038_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X12 c1_n9758_n15640# m3_n9798_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X13 c1_n9758_n15640# m3_n9798_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X14 c1_n9758_n15640# m3_n9798_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X15 c1_n16370_n15640# m3_n16410_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X16 c1_n9758_n15640# m3_n9798_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X17 c1_10078_n15640# m3_10038_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X18 c1_3466_n15640# m3_3426_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X19 c1_n9758_n15640# m3_n9798_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X20 c1_10078_n15640# m3_10038_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X21 c1_n3146_n15640# m3_n3186_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X22 c1_10078_n15640# m3_10038_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X23 c1_n16370_n15640# m3_n16410_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X24 c1_n3146_n15640# m3_n3186_n15680# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
.ends

.subckt sky130_fd_pr__nfet_01v8_4BNSKG a_18_n42# a_n33_n130# a_n76_n42# a_n178_n216#
X0 a_18_n42# a_n33_n130# a_n76_n42# a_n178_n216# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.18
.ends

.subckt sky130_fd_pr__pfet_01v8_X4438S a_18_n72# w_n214_n291# a_n33_n169# a_n76_n72#
X0 a_18_n72# a_n33_n169# a_n76_n72# w_n214_n291# sky130_fd_pr__pfet_01v8 ad=0.2088 pd=2.02 as=0.2088 ps=2.02 w=0.72 l=0.18
.ends

.subckt cs_inv Vp out in Vn VDD VSUBS
XXM1 m1_879_n1632# in out VSUBS sky130_fd_pr__nfet_01v8_4BNSKG
XXM2 m1_917_n552# VDD Vp VDD sky130_fd_pr__pfet_01v8_X4438S
XXM3 out VDD in m1_917_n552# sky130_fd_pr__pfet_01v8_X4438S
XXM4 VSUBS Vn m1_879_n1632# VSUBS sky130_fd_pr__nfet_01v8_4BNSKG
.ends

.subckt sky130_fd_pr__pfet_01v8_HBKBCU w_n214_n399# a_n33_n277# a_n76_n180# a_18_n180#
X0 a_18_n180# a_n33_n277# a_n76_n180# w_n214_n399# sky130_fd_pr__pfet_01v8 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=0.18
.ends

.subckt vco osc vctrl VDD GND
XXM23 GND x1/in osc GND sky130_fd_pr__nfet_01v8_4BNSKG
XXM24 osc VDD x1/in VDD sky130_fd_pr__pfet_01v8_X4438S
Xx1 Vp x7/in x1/in vctrl VDD GND cs_inv
Xx3 Vp x6/in x3/in vctrl VDD GND cs_inv
Xx2 Vp x5/in x2/in vctrl VDD GND cs_inv
Xx4 Vp x3/in x4/in vctrl VDD GND cs_inv
Xx5 Vp x4/in x5/in vctrl VDD GND cs_inv
Xx6 Vp x1/in x6/in vctrl VDD GND cs_inv
Xx7 Vp x2/in x7/in vctrl VDD GND cs_inv
Xsky130_fd_pr__pfet_01v8_HBKBCU_0 VDD Vp VDD Vp sky130_fd_pr__pfet_01v8_HBKBCU
XXM21 GND vctrl Vp GND sky130_fd_pr__nfet_01v8_6FB46G
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_Z926RQ c1_n19676_n37760# c1_n39512_n37760# m3_33180_n37800#
+ m3_n26328_n37800# m3_19956_n37800# c1_n6452_n37760# m3_n6492_n37800# c1_n13064_n37760#
+ m3_6732_n37800# m3_n39552_n37800# m3_13344_n37800# c1_26608_n37760# c1_160_n37760#
+ m3_n19716_n37800# c1_19996_n37760# c1_n32900_n37760# c1_n26288_n37760# m3_120_n37800#
+ c1_33220_n37760# m3_n13104_n37800# c1_13384_n37760# m3_26568_n37800# c1_6772_n37760#
+ m3_n32940_n37800#
X0 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X1 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X2 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X3 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X4 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X5 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X6 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X7 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X8 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X9 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X10 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X11 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X12 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X13 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X14 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X15 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X16 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X17 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X18 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X19 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X20 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X21 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X22 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X23 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X24 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X25 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X26 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X27 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X28 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X29 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X30 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X31 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X32 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X33 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X34 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X35 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X36 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X37 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X38 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X39 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X40 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X41 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X42 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X43 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X44 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X45 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X46 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X47 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X48 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X49 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X50 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X51 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X52 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X53 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X54 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X55 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X56 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X57 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X58 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X59 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X60 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X61 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X62 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X63 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X64 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X65 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X66 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X67 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X68 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X69 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X70 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X71 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X72 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X73 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X74 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X75 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X76 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X77 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X78 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X79 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X80 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X81 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X82 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X83 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X84 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X85 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X86 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X87 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X88 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X89 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X90 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X91 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X92 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X93 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X94 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X95 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X96 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X97 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X98 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X99 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X100 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X101 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X102 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X103 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X104 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X105 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X106 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X107 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X108 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X109 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X110 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X111 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X112 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X113 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X114 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X115 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X116 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X117 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X118 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X119 c1_n39512_n37760# m3_n39552_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X120 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X121 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X122 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X123 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X124 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X125 c1_n26288_n37760# m3_n26328_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X126 c1_6772_n37760# m3_6732_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X127 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X128 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X129 c1_160_n37760# m3_120_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X130 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X131 c1_n19676_n37760# m3_n19716_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X132 c1_26608_n37760# m3_26568_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X133 c1_n32900_n37760# m3_n32940_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X134 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X135 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X136 c1_n13064_n37760# m3_n13104_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X137 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X138 c1_33220_n37760# m3_33180_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X139 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X140 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X141 c1_13384_n37760# m3_13344_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X142 c1_19996_n37760# m3_19956_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X143 c1_n6452_n37760# m3_n6492_n37800# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
.ends

.subckt sky130_fd_pr__pfet_01v8_K9S5FM a_18_n54# w_n214_n273# a_n76_n54# a_n33_n151#
X0 a_18_n54# a_n33_n151# a_n76_n54# w_n214_n273# sky130_fd_pr__pfet_01v8 ad=0.1566 pd=1.66 as=0.1566 ps=1.66 w=0.54 l=0.18
.ends

.subckt cp up vctrl VDD down fd_8_0/VDD fd_8_0/f_out vco_0/VDD fd_8_0/k up_bar2 vco_0/osc
+ vco_0/vctrl down_carry down_b2 GND
XXM12 down_b VDD VDD down sky130_fd_pr__pfet_01v8_KZR7FM
Xsky130_fd_pr__pfet_01v8_K9S7EM_0 up_bar up_bar2 up_bar2 VDD sky130_fd_pr__pfet_01v8_K9S7EM
Xsky130_fd_pr__pfet_01v8_K9S7EM_1 down_b down_b2 down_b2 VDD sky130_fd_pr__pfet_01v8_K9S7EM
XXM18 VDD VDD GND GND sky130_fd_pr__nfet_01v8_6FB46G
XXR2 m1_11512_8746# vctrl sky130_fd_pr__res_generic_po_447X6E
Xfd_8_0 fd_8_0/VDD fd_8_0/k fd_8_0/f_out GND fd_8
XXM3 down_carry down GND GND sky130_fd_pr__nfet_01v8_HAAXKC
XXM4 VDD VDD up_carry up_bar2 sky130_fd_pr__pfet_01v8_7PMXFU
Xsky130_fd_pr__nfet_01v8_6FB27G_0 down_carry down_b2 down_carry down_carry sky130_fd_pr__nfet_01v8_6FB27G
Xsky130_fd_pr__nfet_01v8_6FB46G_0 GND up up_bar GND sky130_fd_pr__nfet_01v8_6FB46G
XXM7 vctrl up_carry up_carry GND sky130_fd_pr__pfet_01v8_KXJ7FM
Xsky130_fd_pr__nfet_01v8_6FB46G_1 down_carry VDD vctrl down_carry sky130_fd_pr__nfet_01v8_6FB46G
Xsky130_fd_pr__nfet_01v8_6FB46G_2 up_bar2 GND up_bar up_bar2 sky130_fd_pr__nfet_01v8_6FB46G
Xsky130_fd_pr__cap_mim_m3_1_39XMLG_0 GND vctrl vctrl vctrl vctrl GND GND vctrl GND
+ GND sky130_fd_pr__cap_mim_m3_1_39XMLG
Xsky130_fd_pr__nfet_01v8_6FB46G_3 GND down down_b GND sky130_fd_pr__nfet_01v8_6FB46G
Xsky130_fd_pr__nfet_01v8_6FB46G_5 down_b2 GND down_b down_b2 sky130_fd_pr__nfet_01v8_6FB46G
Xsky130_fd_pr__pfet_01v8_KZR7FM_0 VDD VDD GND GND sky130_fd_pr__pfet_01v8_KZR7FM
Xsky130_fd_pr__pfet_01v8_KZR7FM_1 up_bar VDD VDD up sky130_fd_pr__pfet_01v8_KZR7FM
Xvco_0 vco_0/osc vco_0/vctrl vco_0/VDD GND vco
Xsky130_fd_pr__cap_mim_m3_1_Z926RQ_0 m1_11512_8746# m1_11512_8746# GND GND GND m1_11512_8746#
+ GND m1_11512_8746# GND GND GND m1_11512_8746# m1_11512_8746# GND m1_11512_8746#
+ m1_11512_8746# m1_11512_8746# GND m1_11512_8746# GND m1_11512_8746# GND m1_11512_8746#
+ GND sky130_fd_pr__cap_mim_m3_1_Z926RQ
XXM10 up_carry up_carry up_carry up sky130_fd_pr__pfet_01v8_K9S5FM
.ends

.subckt pll VDD GND f_clk_in f_clk_out
Xpfd_lay_0 f_clk_in VDD pfd_lay_0/f_vco cp_0/down cp_0/up GND pfd_lay
Xcp_0 cp_0/up cp_0/vctrl VDD cp_0/down VDD pfd_lay_0/f_vco VDD f_clk_out cp_0/up_bar2
+ f_clk_out cp_0/vctrl cp_0/down_carry cp_0/down_b2 GND cp
.ends

