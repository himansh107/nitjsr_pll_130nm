magic
tech sky130A
magscale 1 2
timestamp 1714832304
<< nwell >>
rect 1556 581 5094 902
rect 1885 -132 2260 -131
rect 2514 -132 2716 -131
rect 1885 -452 2716 -132
rect 4195 -581 4688 -260
rect 1503 -2003 5388 -1682
rect 2147 -2924 2910 -2603
<< locali >>
rect 2635 744 2785 746
rect 2635 696 2636 744
rect 2684 696 2785 744
rect 2635 695 2785 696
rect 2740 580 2778 695
rect 1230 540 1440 580
rect 1490 540 2140 580
rect 2260 577 2470 580
rect 2260 543 2433 577
rect 2467 543 2470 577
rect 2260 540 2470 543
rect 2740 540 3010 580
rect 3060 540 3660 580
rect 3980 570 4020 720
rect 4920 650 5010 690
rect 4970 580 5010 650
rect 2740 440 2780 540
rect 3700 530 4020 570
rect 4150 530 4330 570
rect 2200 400 2780 440
rect 4150 397 4190 530
rect 4560 530 4820 580
rect 4970 540 5210 580
rect 5270 540 5540 580
rect 5580 540 5590 580
rect 4771 520 4810 530
rect 4970 430 5010 540
rect 4150 363 4153 397
rect 4187 363 4190 397
rect 4480 390 5010 430
rect 4150 360 4190 363
rect 2070 10 2310 50
rect 2830 0 3140 40
rect 1680 -93 1960 -90
rect 1680 -127 1683 -93
rect 1717 -127 1960 -93
rect 1680 -130 1960 -127
rect 2100 -130 2430 -90
rect 2570 -120 2740 -80
rect 2883 -117 3003 -83
rect 2285 -150 2325 -130
rect 2285 -190 2288 -150
rect 2322 -190 2325 -150
rect 3720 -323 3760 -320
rect 3720 -357 3723 -323
rect 3757 -357 3760 -323
rect 3720 -450 3760 -357
rect 3720 -490 3870 -450
rect 3528 -590 3952 -588
rect 3528 -593 4100 -590
rect 4420 -593 4970 -590
rect 3528 -627 3533 -593
rect 3567 -627 4100 -593
rect 4420 -627 4933 -593
rect 4967 -627 4970 -593
rect 3528 -630 4100 -627
rect 4420 -630 4970 -627
rect 3528 -632 3952 -630
rect 3740 -760 3920 -720
rect 3741 -993 3779 -760
rect 3741 -1027 3743 -993
rect 3777 -1027 3779 -993
rect 3741 -1029 3779 -1027
rect 1420 -2040 1634 -2000
rect 2450 -2003 2650 -2000
rect 1680 -2050 2330 -2010
rect 2450 -2037 2613 -2003
rect 2647 -2037 2650 -2003
rect 2450 -2040 2650 -2037
rect 2970 -2040 3190 -2000
rect 3240 -2040 3830 -2000
rect 2840 -2053 2880 -2050
rect 2840 -2087 2843 -2053
rect 2877 -2087 2880 -2053
rect 2840 -2140 2880 -2087
rect 2970 -2140 3010 -2040
rect 3920 -2050 4250 -2010
rect 4290 -2050 4300 -2010
rect 4340 -2013 4520 -2010
rect 4340 -2047 4343 -2013
rect 4377 -2047 4520 -2013
rect 4340 -2050 4520 -2047
rect 4753 -2047 4922 -2013
rect 5140 -2013 5270 -2010
rect 5140 -2047 5387 -2013
rect 5140 -2050 5270 -2047
rect 5450 -2050 5940 -2010
rect 2420 -2180 3010 -2140
rect 5230 -2150 5270 -2050
rect 4650 -2190 5270 -2150
rect 2000 -2510 2270 -2470
rect 2470 -2480 2870 -2440
rect 2470 -2560 2510 -2480
rect 1947 -2607 2237 -2573
rect 2360 -2600 2510 -2560
rect 2580 -2700 2620 -2480
rect 2747 -2607 2857 -2573
rect 3000 -2610 3300 -2570
<< viali >>
rect 2636 696 2684 744
rect 3980 720 4020 760
rect 1190 540 1230 580
rect 2433 543 2467 577
rect 4880 650 4920 690
rect 4453 523 4487 557
rect 5540 540 5580 580
rect 4771 481 4810 520
rect 4153 363 4187 397
rect 2310 10 2350 50
rect 3140 0 3180 40
rect 1683 -127 1717 -93
rect 2430 -130 2470 -90
rect 2530 -120 2570 -80
rect 3003 -117 3037 -83
rect 2288 -190 2322 -150
rect 3723 -357 3757 -323
rect 3870 -490 3910 -450
rect 3533 -627 3567 -593
rect 4153 -627 4187 -593
rect 4933 -627 4967 -593
rect 3920 -760 3960 -720
rect 4233 -757 4267 -723
rect 4354 -735 4388 -701
rect 3743 -1027 3777 -993
rect 1380 -2040 1420 -2000
rect 2613 -2037 2647 -2003
rect 2843 -2087 2877 -2053
rect 4250 -2050 4290 -2010
rect 4343 -2047 4377 -2013
rect 4653 -2057 4687 -2023
rect 4922 -2047 4956 -2013
rect 5100 -2050 5140 -2010
rect 5940 -2050 5980 -2010
rect 1960 -2510 2000 -2470
rect 1913 -2607 1947 -2573
rect 2713 -2607 2747 -2573
rect 3300 -2610 3340 -2570
rect 2580 -2740 2620 -2700
<< metal1 >>
rect 2424 1316 2476 1322
rect 4868 1310 4874 1316
rect 2476 1270 4874 1310
rect 4868 1264 4874 1270
rect 4926 1264 4932 1316
rect 2424 1258 2476 1264
rect 3312 1048 3512 1220
rect 6946 1140 6998 1146
rect 6690 1134 6696 1140
rect 6560 1094 6696 1134
rect 1380 952 5408 1048
rect 1380 884 5520 952
rect 4874 826 4926 832
rect 2418 724 2424 776
rect 2476 724 2482 776
rect 4874 768 4926 774
rect 3968 760 4032 766
rect 2630 744 2690 756
rect 850 580 1050 676
rect 1184 580 1236 592
rect 2430 583 2470 724
rect 2630 696 2636 744
rect 2684 696 2690 744
rect 3968 720 3980 760
rect 4020 720 4490 760
rect 3968 714 4032 720
rect 2630 620 2690 696
rect 850 540 1190 580
rect 1230 540 1236 580
rect 850 476 1050 540
rect 1184 528 1236 540
rect 2421 577 2479 583
rect 2421 543 2433 577
rect 2467 543 2479 577
rect 2624 560 2630 620
rect 2690 560 2696 620
rect 4450 569 4490 720
rect 4880 702 4920 768
rect 4874 690 4926 702
rect 4874 650 4880 690
rect 4920 650 4926 690
rect 4874 638 4926 650
rect 5534 580 5586 592
rect 6560 580 6600 1094
rect 6690 1088 6696 1094
rect 6748 1088 6754 1140
rect 6998 1094 7172 1134
rect 6946 1082 6998 1088
rect 2421 537 2479 543
rect 4447 557 4493 569
rect 4447 523 4453 557
rect 4487 523 4493 557
rect 5534 540 5540 580
rect 5580 540 6600 580
rect 4765 527 4817 533
rect 5534 528 5586 540
rect 4447 511 4493 523
rect 4759 475 4765 526
rect 4817 475 4822 526
rect 4765 469 4817 475
rect 3928 354 3934 406
rect 3986 400 3992 406
rect 4141 400 4199 403
rect 3986 397 4199 400
rect 3986 363 4153 397
rect 4187 363 4199 397
rect 3986 360 4199 363
rect 3986 354 3992 360
rect 4141 357 4199 360
rect 1380 272 5408 300
rect 1380 204 5520 272
rect 1380 136 5408 204
rect 2304 56 2356 62
rect 2304 -2 2356 4
rect 2424 56 2476 62
rect 2988 34 2994 86
rect 3046 34 3052 86
rect 3134 40 3186 52
rect 2424 -2 2476 4
rect 2430 -78 2470 -2
rect 1671 -93 1729 -87
rect 1671 -127 1683 -93
rect 1717 -127 1729 -93
rect 1671 -133 1729 -127
rect 2424 -90 2476 -78
rect 2424 -130 2430 -90
rect 2470 -130 2476 -90
rect 1680 -710 1720 -133
rect 2282 -144 2334 -138
rect 2424 -142 2476 -130
rect 2524 -80 2576 -68
rect 3004 -71 3036 34
rect 3134 0 3140 40
rect 3180 0 3186 40
rect 3404 0 3604 136
rect 3928 34 3934 86
rect 3986 34 3992 86
rect 3134 -12 3186 0
rect 2524 -120 2530 -80
rect 2570 -120 2576 -80
rect 2524 -132 2576 -120
rect 2997 -83 3043 -71
rect 2997 -117 3003 -83
rect 3037 -117 3043 -83
rect 2997 -129 3043 -117
rect 2276 -196 2282 -144
rect 2282 -202 2334 -196
rect 2289 -375 2295 -323
rect 2347 -331 2353 -323
rect 2532 -331 2569 -132
rect 2347 -368 2569 -331
rect 2347 -375 2353 -368
rect 1840 -544 3036 -408
rect 2484 -680 2684 -544
rect 3140 -710 3180 -12
rect 3940 -30 3980 34
rect 3940 -70 4970 -30
rect 3714 -144 3766 -138
rect 3714 -202 3766 -196
rect 3720 -311 3760 -202
rect 4160 -300 4360 -100
rect 3717 -323 3763 -311
rect 3717 -357 3723 -323
rect 3757 -357 3763 -323
rect 4450 -350 4644 -250
rect 3717 -369 3763 -357
rect 3864 -450 3916 -438
rect 3864 -490 3870 -450
rect 3910 -490 4190 -450
rect 3864 -502 3916 -490
rect 4150 -581 4190 -490
rect 4930 -581 4970 -70
rect 3521 -593 3579 -587
rect 3521 -627 3533 -593
rect 3567 -627 3579 -593
rect 3521 -633 3579 -627
rect 4147 -593 4193 -581
rect 4147 -627 4153 -593
rect 4187 -627 4193 -593
rect 1680 -750 3180 -710
rect 2290 -855 2296 -803
rect 2348 -855 2354 -803
rect 2304 -1109 2341 -855
rect 2728 -1006 2734 -954
rect 2786 -958 2792 -954
rect 3528 -958 3572 -633
rect 4147 -639 4193 -627
rect 4927 -593 4973 -581
rect 4927 -627 4933 -593
rect 4967 -627 4973 -593
rect 4927 -639 4973 -627
rect 4485 -693 4537 -687
rect 4342 -700 4400 -695
rect 4342 -701 4485 -700
rect 3914 -720 3966 -708
rect 4221 -720 4279 -717
rect 3914 -760 3920 -720
rect 3960 -723 4279 -720
rect 3960 -757 4233 -723
rect 4267 -757 4279 -723
rect 4342 -735 4354 -701
rect 4388 -735 4485 -701
rect 4342 -737 4485 -735
rect 4342 -741 4400 -737
rect 4485 -751 4537 -745
rect 3960 -760 4279 -757
rect 3914 -772 3966 -760
rect 4221 -763 4279 -760
rect 4450 -850 4644 -790
rect 2786 -1002 3572 -958
rect 4270 -890 4644 -850
rect 3731 -991 3789 -987
rect 4128 -991 4134 -984
rect 3731 -993 4134 -991
rect 2786 -1006 2792 -1002
rect 3731 -1027 3743 -993
rect 3777 -1027 4134 -993
rect 3731 -1029 4134 -1027
rect 3731 -1033 3789 -1029
rect 4128 -1036 4134 -1029
rect 4186 -1036 4192 -984
rect 4270 -1050 4470 -890
rect 4628 -1109 4634 -1101
rect 2304 -1146 4634 -1109
rect 2304 -1481 2341 -1146
rect 4628 -1153 4634 -1146
rect 4686 -1153 4692 -1101
rect 1132 -1518 2341 -1481
rect 2610 -1320 5140 -1280
rect 2610 -1498 2650 -1320
rect 2604 -1504 2656 -1498
rect 650 -2000 850 -1940
rect 964 -1994 1016 -1988
rect 650 -2040 964 -2000
rect 650 -2140 850 -2040
rect 964 -2052 1016 -2046
rect 1133 -2914 1167 -1518
rect 2604 -1562 2656 -1556
rect 3588 -1605 3788 -1432
rect 5100 -1494 5140 -1320
rect 5088 -1546 5094 -1494
rect 5146 -1546 5152 -1494
rect 1566 -1632 5594 -1605
rect 1566 -1700 5704 -1632
rect 1566 -1769 5630 -1700
rect 5580 -1770 5630 -1769
rect 5094 -1804 5146 -1798
rect 2598 -1866 2604 -1814
rect 2656 -1866 2662 -1814
rect 4250 -1850 4690 -1810
rect 2834 -1858 2886 -1852
rect 1238 -2046 1244 -1994
rect 1296 -2000 1302 -1994
rect 1374 -2000 1426 -1988
rect 2610 -1997 2650 -1866
rect 2834 -1916 2886 -1910
rect 1296 -2040 1380 -2000
rect 1420 -2040 1426 -2000
rect 1296 -2046 1302 -2040
rect 1374 -2052 1426 -2040
rect 2601 -2003 2659 -1997
rect 2601 -2037 2613 -2003
rect 2647 -2037 2659 -2003
rect 2728 -2006 2734 -1954
rect 2786 -1960 2792 -1954
rect 2840 -1960 2880 -1916
rect 2786 -2000 2880 -1960
rect 2786 -2006 2792 -2000
rect 2601 -2043 2659 -2037
rect 2840 -2047 2880 -2000
rect 4250 -2004 4290 -1850
rect 4238 -2010 4302 -2004
rect 2831 -2053 2889 -2047
rect 2831 -2087 2843 -2053
rect 2877 -2087 2889 -2053
rect 4238 -2050 4250 -2010
rect 4290 -2050 4302 -2010
rect 4238 -2056 4302 -2050
rect 4331 -2013 4389 -2007
rect 4650 -2011 4690 -1850
rect 4907 -1866 4913 -1814
rect 4965 -1866 4971 -1814
rect 5094 -1862 5146 -1856
rect 4922 -2001 4956 -1866
rect 5100 -1998 5140 -1862
rect 4331 -2047 4343 -2013
rect 4377 -2047 4389 -2013
rect 4331 -2053 4389 -2047
rect 4647 -2023 4693 -2011
rect 2831 -2093 2889 -2087
rect 4340 -2124 4380 -2053
rect 4647 -2057 4653 -2023
rect 4687 -2057 4693 -2023
rect 4647 -2069 4693 -2057
rect 4916 -2013 4962 -2001
rect 4916 -2047 4922 -2013
rect 4956 -2047 4962 -2013
rect 4916 -2059 4962 -2047
rect 5094 -2010 5146 -1998
rect 5094 -2050 5100 -2010
rect 5140 -2050 5146 -2010
rect 5094 -2062 5146 -2050
rect 5934 -2010 5986 -1998
rect 7306 -2004 7358 -1998
rect 7034 -2010 7040 -2004
rect 5934 -2050 5940 -2010
rect 5980 -2050 7040 -2010
rect 5934 -2062 5986 -2050
rect 7034 -2056 7040 -2050
rect 7092 -2056 7098 -2004
rect 7410 -2010 7450 -1632
rect 7358 -2050 7450 -2010
rect 7306 -2062 7358 -2056
rect 4328 -2176 4334 -2124
rect 4386 -2176 4392 -2124
rect 5580 -2216 5640 -2210
rect 1622 -2244 5640 -2216
rect 1472 -2312 5704 -2244
rect 1472 -2380 5602 -2312
rect 3294 -2424 3346 -2418
rect 1954 -2464 2006 -2458
rect 2698 -2496 2704 -2444
rect 2756 -2496 2762 -2444
rect 3294 -2482 3346 -2476
rect 4134 -2434 4186 -2428
rect 1954 -2522 2006 -2516
rect 2713 -2561 2747 -2496
rect 1901 -2573 1959 -2567
rect 1901 -2607 1913 -2573
rect 1947 -2607 1959 -2573
rect 1901 -2613 1959 -2607
rect 2707 -2573 2753 -2561
rect 3300 -2564 3340 -2482
rect 4134 -2492 4186 -2486
rect 4334 -2454 4386 -2448
rect 2707 -2607 2713 -2573
rect 2747 -2607 2753 -2573
rect 1914 -2914 1946 -2613
rect 2707 -2619 2753 -2607
rect 3288 -2570 3352 -2564
rect 3288 -2610 3300 -2570
rect 3340 -2610 3352 -2570
rect 3288 -2616 3352 -2610
rect 2568 -2700 2632 -2694
rect 4140 -2700 4180 -2492
rect 5000 -2480 5200 -2380
rect 4334 -2512 4386 -2506
rect 4340 -2700 4380 -2512
rect 2568 -2740 2580 -2700
rect 2620 -2740 4380 -2700
rect 2568 -2746 2632 -2740
rect 1133 -2946 1946 -2914
rect 1133 -2947 1167 -2946
rect 2116 -2992 3128 -2924
rect 2668 -3176 2868 -2992
<< via1 >>
rect 2424 1264 2476 1316
rect 4874 1264 4926 1316
rect 2424 724 2476 776
rect 4874 774 4926 826
rect 2630 560 2690 620
rect 6696 1088 6748 1140
rect 6946 1088 6998 1140
rect 4765 520 4817 527
rect 4765 481 4771 520
rect 4771 481 4810 520
rect 4810 481 4817 520
rect 4765 475 4817 481
rect 3934 354 3986 406
rect 2304 50 2356 56
rect 2304 10 2310 50
rect 2310 10 2350 50
rect 2350 10 2356 50
rect 2304 4 2356 10
rect 2424 4 2476 56
rect 2994 34 3046 86
rect 3934 34 3986 86
rect 2282 -150 2334 -144
rect 2282 -190 2288 -150
rect 2288 -190 2322 -150
rect 2322 -190 2334 -150
rect 2282 -196 2334 -190
rect 2295 -375 2347 -323
rect 3714 -196 3766 -144
rect 2296 -855 2348 -803
rect 2734 -1006 2786 -954
rect 4485 -745 4537 -693
rect 4134 -1036 4186 -984
rect 4634 -1153 4686 -1101
rect 964 -2046 1016 -1994
rect 2604 -1556 2656 -1504
rect 5094 -1546 5146 -1494
rect 2604 -1866 2656 -1814
rect 1244 -2046 1296 -1994
rect 2834 -1910 2886 -1858
rect 2734 -2006 2786 -1954
rect 4913 -1866 4965 -1814
rect 5094 -1856 5146 -1804
rect 7040 -2056 7092 -2004
rect 7306 -2056 7358 -2004
rect 4334 -2176 4386 -2124
rect 1954 -2470 2006 -2464
rect 1954 -2510 1960 -2470
rect 1960 -2510 2000 -2470
rect 2000 -2510 2006 -2470
rect 2704 -2496 2756 -2444
rect 3294 -2476 3346 -2424
rect 1954 -2516 2006 -2510
rect 4134 -2486 4186 -2434
rect 4334 -2506 4386 -2454
<< metal2 >>
rect 4874 1316 4926 1322
rect 2418 1264 2424 1316
rect 2476 1264 2482 1316
rect 2430 782 2470 1264
rect 4874 1258 4926 1264
rect 4880 826 4920 1258
rect 6696 1140 6748 1146
rect 6940 1134 6946 1140
rect 6748 1094 6946 1134
rect 6940 1088 6946 1094
rect 6998 1088 7004 1140
rect 6696 1082 6748 1088
rect 2424 776 2476 782
rect 4868 774 4874 826
rect 4926 774 4932 826
rect 2424 718 2476 724
rect 2630 620 2690 626
rect 2422 370 2478 377
rect 2630 370 2690 560
rect 4759 475 4765 527
rect 4817 475 4823 527
rect 2420 368 2690 370
rect 2420 312 2422 368
rect 2478 312 2690 368
rect 3934 406 3986 412
rect 3934 348 3986 354
rect 2420 310 2690 312
rect 2422 303 2478 310
rect 3940 240 3980 348
rect 2310 200 3980 240
rect 2310 56 2350 200
rect 3000 92 3040 200
rect 3940 92 3980 200
rect 2994 86 3046 92
rect 2420 60 2480 69
rect 2298 4 2304 56
rect 2356 4 2362 56
rect 2418 4 2420 56
rect 2480 4 2482 56
rect 2994 28 3046 34
rect 3934 86 3986 92
rect 3934 28 3986 34
rect 2420 -9 2480 0
rect 4772 -99 4811 475
rect 2276 -196 2282 -144
rect 2334 -150 2340 -144
rect 3708 -150 3714 -144
rect 2334 -190 3714 -150
rect 2334 -196 2340 -190
rect 3708 -196 3714 -190
rect 3766 -196 3772 -144
rect 2295 -323 2347 -317
rect 2295 -381 2347 -375
rect 2303 -797 2340 -381
rect 4479 -745 4485 -693
rect 4537 -701 4543 -693
rect 4773 -701 4810 -99
rect 4537 -738 4810 -701
rect 4537 -745 4543 -738
rect 2296 -803 2348 -797
rect 2296 -861 2348 -855
rect 2734 -954 2786 -948
rect 2734 -1012 2786 -1006
rect 4134 -984 4186 -978
rect 2738 -1472 2782 -1012
rect 4134 -1042 4186 -1036
rect 2598 -1556 2604 -1504
rect 2656 -1556 2662 -1504
rect 2610 -1808 2650 -1556
rect 2604 -1814 2656 -1808
rect 2604 -1872 2656 -1866
rect 2740 -1948 2780 -1472
rect 2828 -1910 2834 -1858
rect 2886 -1864 2892 -1858
rect 2952 -1864 3340 -1860
rect 2886 -1900 3340 -1864
rect 2886 -1904 2982 -1900
rect 2886 -1910 2892 -1904
rect 2734 -1954 2786 -1948
rect 1244 -1994 1296 -1988
rect 958 -2046 964 -1994
rect 1016 -2000 1022 -1994
rect 1016 -2040 1244 -2000
rect 1016 -2046 1022 -2040
rect 2734 -2012 2786 -2006
rect 1244 -2052 1296 -2046
rect 1960 -2300 2750 -2260
rect 1960 -2464 2000 -2300
rect 2710 -2438 2750 -2300
rect 3300 -2424 3340 -1900
rect 2704 -2444 2756 -2438
rect 1948 -2516 1954 -2464
rect 2006 -2516 2012 -2464
rect 3288 -2476 3294 -2424
rect 3346 -2476 3352 -2424
rect 4140 -2434 4180 -1042
rect 4634 -1101 4686 -1095
rect 4773 -1108 4810 -738
rect 4686 -1145 4810 -1108
rect 4634 -1159 4686 -1153
rect 4773 -1461 4810 -1145
rect 4773 -1498 4958 -1461
rect 5094 -1494 5146 -1488
rect 4922 -1808 4956 -1498
rect 5094 -1552 5146 -1546
rect 5100 -1804 5140 -1552
rect 4913 -1814 4965 -1808
rect 5088 -1856 5094 -1804
rect 5146 -1856 5152 -1804
rect 4913 -1872 4965 -1866
rect 7040 -2004 7092 -1998
rect 7300 -2010 7306 -2004
rect 7092 -2050 7306 -2010
rect 7300 -2056 7306 -2050
rect 7358 -2056 7364 -2004
rect 7040 -2062 7092 -2056
rect 4334 -2124 4386 -2118
rect 4334 -2182 4386 -2176
rect 4128 -2486 4134 -2434
rect 4186 -2486 4192 -2434
rect 4340 -2454 4380 -2182
rect 2704 -2502 2756 -2496
rect 4328 -2506 4334 -2454
rect 4386 -2506 4392 -2454
<< via2 >>
rect 2422 312 2478 368
rect 2420 56 2480 60
rect 2420 4 2424 56
rect 2424 4 2476 56
rect 2476 4 2480 56
rect 2420 0 2480 4
<< metal3 >>
rect 2417 368 2483 373
rect 2417 312 2422 368
rect 2478 312 2483 368
rect 2417 307 2483 312
rect 2420 65 2480 307
rect 2415 60 2485 65
rect 2415 0 2420 60
rect 2480 0 2485 60
rect 2415 -5 2485 0
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 3534 0 1 320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1709947739
transform 1 0 2890 0 1 320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1709947739
transform 1 0 1326 0 1 320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1709947739
transform 1 0 5098 0 1 320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 2062 0 1 320
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 4270 0 1 320
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 4602 0 1 -842
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1709947739
transform 1 0 5616 0 1 -2262
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1709947739
transform 1 0 1764 0 -1 126
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1709947739
transform 1 0 3118 0 -1 -2368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1709947739
transform 1 0 5374 0 1 320
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1709947739
transform 1 0 4018 0 1 -842
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  x2
timestamp 1709947739
transform -1 0 2430 0 -1 -2342
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1709947739
transform 1 0 1510 0 1 -2264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  x5
timestamp 1709947739
transform 1 0 4454 0 1 -2264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  x6
timestamp 1709947739
transform 1 0 2246 0 1 -2264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x8
timestamp 1709947739
transform 1 0 1892 0 -1 130
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x9
timestamp 1709947739
transform 1 0 2662 0 -1 140
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x10
timestamp 1709947739
transform 1 0 3074 0 1 -2264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  x11
timestamp 1709947739
transform -1 0 3076 0 -1 -2354
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x12
timestamp 1709947739
transform 1 0 3718 0 1 -2264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x13
timestamp 1709947739
transform 1 0 5282 0 1 -2264
box -38 -48 314 592
<< labels >>
flabel metal1 850 476 1050 676 0 FreeSans 256 0 0 0 f_clk_in
port 0 nsew
flabel metal1 5000 -2480 5200 -2280 0 FreeSans 256 0 0 0 VGND
port 3 nsew
flabel metal1 4270 -1050 4470 -850 0 FreeSans 256 0 0 0 VGND
port 3 nsew
flabel metal1 3404 0 3604 200 0 FreeSans 256 0 0 0 VGND
port 3 nsew
flabel metal1 2484 -680 2684 -480 0 FreeSans 256 0 0 0 VPWR
port 2 nsew
flabel metal1 3588 -1632 3788 -1432 0 FreeSans 256 0 0 0 VPWR
port 2 nsew
flabel metal1 2668 -3176 2868 -2976 0 FreeSans 256 0 0 0 VPWR
port 2 nsew
flabel metal1 4160 -300 4360 -100 0 FreeSans 256 0 0 0 VPWR
port 2 nsew
flabel metal1 3312 1020 3512 1220 0 FreeSans 256 0 0 0 VPWR
port 2 nsew
flabel metal1 s 2088 916 2122 950 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 2060 885 2336 981 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 2917 916 2951 950 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 2888 885 3164 981 1 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 3561 916 3595 950 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 3532 885 3808 981 1 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 4298 916 4332 950 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 4268 885 4636 981 1 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 5125 916 5159 950 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 5096 885 5372 981 1 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 650 -2140 850 -1940 0 FreeSans 256 0 0 0 f_vco
port 5 nsew
flabel locali 1692 554 1692 554 0 FreeSans 256 0 0 0 test1
flabel locali 2502 418 2502 418 0 FreeSans 256 0 0 0 test2
flabel space 2908 1290 2908 1290 0 FreeSans 256 0 0 0 test3
flabel locali 3866 546 3866 546 0 FreeSans 256 0 0 0 test4
<< end >>
