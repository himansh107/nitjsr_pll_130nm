VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__cap_mim_m3_1_Z926RQ
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_mim_m3_1_Z926RQ ;
  ORIGIN -165.900 -158.600 ;
  SIZE 30.400 BY 30.400 ;
  OBS
      LAYER met3 ;
        RECT -197.760 158.600 -165.900 189.000 ;
        RECT -164.700 158.600 -132.840 189.000 ;
        RECT -131.640 158.600 -99.780 189.000 ;
        RECT -98.580 158.600 -66.720 189.000 ;
        RECT -65.520 158.600 -33.660 189.000 ;
        RECT -32.460 158.600 -0.600 189.000 ;
        RECT 0.600 158.600 32.460 189.000 ;
        RECT 33.660 158.600 65.520 189.000 ;
        RECT 66.720 158.600 98.580 189.000 ;
        RECT 99.780 158.600 131.640 189.000 ;
        RECT 132.840 158.600 164.700 189.000 ;
        RECT 165.900 158.600 197.760 189.000 ;
        RECT -197.760 127.000 -165.900 157.400 ;
        RECT -164.700 127.000 -132.840 157.400 ;
        RECT -131.640 127.000 -99.780 157.400 ;
        RECT -98.580 127.000 -66.720 157.400 ;
        RECT -65.520 127.000 -33.660 157.400 ;
        RECT -32.460 127.000 -0.600 157.400 ;
        RECT 0.600 127.000 32.460 157.400 ;
        RECT 33.660 127.000 65.520 157.400 ;
        RECT 66.720 127.000 98.580 157.400 ;
        RECT 99.780 127.000 131.640 157.400 ;
        RECT 132.840 127.000 164.700 157.400 ;
        RECT 165.900 127.000 197.760 157.400 ;
        RECT -197.760 95.400 -165.900 125.800 ;
        RECT -164.700 95.400 -132.840 125.800 ;
        RECT -131.640 95.400 -99.780 125.800 ;
        RECT -98.580 95.400 -66.720 125.800 ;
        RECT -65.520 95.400 -33.660 125.800 ;
        RECT -32.460 95.400 -0.600 125.800 ;
        RECT 0.600 95.400 32.460 125.800 ;
        RECT 33.660 95.400 65.520 125.800 ;
        RECT 66.720 95.400 98.580 125.800 ;
        RECT 99.780 95.400 131.640 125.800 ;
        RECT 132.840 95.400 164.700 125.800 ;
        RECT 165.900 95.400 197.760 125.800 ;
        RECT -197.760 63.800 -165.900 94.200 ;
        RECT -164.700 63.800 -132.840 94.200 ;
        RECT -131.640 63.800 -99.780 94.200 ;
        RECT -98.580 63.800 -66.720 94.200 ;
        RECT -65.520 63.800 -33.660 94.200 ;
        RECT -32.460 63.800 -0.600 94.200 ;
        RECT 0.600 63.800 32.460 94.200 ;
        RECT 33.660 63.800 65.520 94.200 ;
        RECT 66.720 63.800 98.580 94.200 ;
        RECT 99.780 63.800 131.640 94.200 ;
        RECT 132.840 63.800 164.700 94.200 ;
        RECT 165.900 63.800 197.760 94.200 ;
        RECT -197.760 32.200 -165.900 62.600 ;
        RECT -164.700 32.200 -132.840 62.600 ;
        RECT -131.640 32.200 -99.780 62.600 ;
        RECT -98.580 32.200 -66.720 62.600 ;
        RECT -65.520 32.200 -33.660 62.600 ;
        RECT -32.460 32.200 -0.600 62.600 ;
        RECT 0.600 32.200 32.460 62.600 ;
        RECT 33.660 32.200 65.520 62.600 ;
        RECT 66.720 32.200 98.580 62.600 ;
        RECT 99.780 32.200 131.640 62.600 ;
        RECT 132.840 32.200 164.700 62.600 ;
        RECT 165.900 32.200 197.760 62.600 ;
        RECT -197.760 0.600 -165.900 31.000 ;
        RECT -164.700 0.600 -132.840 31.000 ;
        RECT -131.640 0.600 -99.780 31.000 ;
        RECT -98.580 0.600 -66.720 31.000 ;
        RECT -65.520 0.600 -33.660 31.000 ;
        RECT -32.460 0.600 -0.600 31.000 ;
        RECT 0.600 0.600 32.460 31.000 ;
        RECT 33.660 0.600 65.520 31.000 ;
        RECT 66.720 0.600 98.580 31.000 ;
        RECT 99.780 0.600 131.640 31.000 ;
        RECT 132.840 0.600 164.700 31.000 ;
        RECT 165.900 0.600 197.760 31.000 ;
        RECT -197.760 -31.000 -165.900 -0.600 ;
        RECT -164.700 -31.000 -132.840 -0.600 ;
        RECT -131.640 -31.000 -99.780 -0.600 ;
        RECT -98.580 -31.000 -66.720 -0.600 ;
        RECT -65.520 -31.000 -33.660 -0.600 ;
        RECT -32.460 -31.000 -0.600 -0.600 ;
        RECT 0.600 -31.000 32.460 -0.600 ;
        RECT 33.660 -31.000 65.520 -0.600 ;
        RECT 66.720 -31.000 98.580 -0.600 ;
        RECT 99.780 -31.000 131.640 -0.600 ;
        RECT 132.840 -31.000 164.700 -0.600 ;
        RECT 165.900 -31.000 197.760 -0.600 ;
        RECT -197.760 -62.600 -165.900 -32.200 ;
        RECT -164.700 -62.600 -132.840 -32.200 ;
        RECT -131.640 -62.600 -99.780 -32.200 ;
        RECT -98.580 -62.600 -66.720 -32.200 ;
        RECT -65.520 -62.600 -33.660 -32.200 ;
        RECT -32.460 -62.600 -0.600 -32.200 ;
        RECT 0.600 -62.600 32.460 -32.200 ;
        RECT 33.660 -62.600 65.520 -32.200 ;
        RECT 66.720 -62.600 98.580 -32.200 ;
        RECT 99.780 -62.600 131.640 -32.200 ;
        RECT 132.840 -62.600 164.700 -32.200 ;
        RECT 165.900 -62.600 197.760 -32.200 ;
        RECT -197.760 -94.200 -165.900 -63.800 ;
        RECT -164.700 -94.200 -132.840 -63.800 ;
        RECT -131.640 -94.200 -99.780 -63.800 ;
        RECT -98.580 -94.200 -66.720 -63.800 ;
        RECT -65.520 -94.200 -33.660 -63.800 ;
        RECT -32.460 -94.200 -0.600 -63.800 ;
        RECT 0.600 -94.200 32.460 -63.800 ;
        RECT 33.660 -94.200 65.520 -63.800 ;
        RECT 66.720 -94.200 98.580 -63.800 ;
        RECT 99.780 -94.200 131.640 -63.800 ;
        RECT 132.840 -94.200 164.700 -63.800 ;
        RECT 165.900 -94.200 197.760 -63.800 ;
        RECT -197.760 -125.800 -165.900 -95.400 ;
        RECT -164.700 -125.800 -132.840 -95.400 ;
        RECT -131.640 -125.800 -99.780 -95.400 ;
        RECT -98.580 -125.800 -66.720 -95.400 ;
        RECT -65.520 -125.800 -33.660 -95.400 ;
        RECT -32.460 -125.800 -0.600 -95.400 ;
        RECT 0.600 -125.800 32.460 -95.400 ;
        RECT 33.660 -125.800 65.520 -95.400 ;
        RECT 66.720 -125.800 98.580 -95.400 ;
        RECT 99.780 -125.800 131.640 -95.400 ;
        RECT 132.840 -125.800 164.700 -95.400 ;
        RECT 165.900 -125.800 197.760 -95.400 ;
        RECT -197.760 -157.400 -165.900 -127.000 ;
        RECT -164.700 -157.400 -132.840 -127.000 ;
        RECT -131.640 -157.400 -99.780 -127.000 ;
        RECT -98.580 -157.400 -66.720 -127.000 ;
        RECT -65.520 -157.400 -33.660 -127.000 ;
        RECT -32.460 -157.400 -0.600 -127.000 ;
        RECT 0.600 -157.400 32.460 -127.000 ;
        RECT 33.660 -157.400 65.520 -127.000 ;
        RECT 66.720 -157.400 98.580 -127.000 ;
        RECT 99.780 -157.400 131.640 -127.000 ;
        RECT 132.840 -157.400 164.700 -127.000 ;
        RECT 165.900 -157.400 197.760 -127.000 ;
        RECT -197.760 -189.000 -165.900 -158.600 ;
        RECT -164.700 -189.000 -132.840 -158.600 ;
        RECT -131.640 -189.000 -99.780 -158.600 ;
        RECT -98.580 -189.000 -66.720 -158.600 ;
        RECT -65.520 -189.000 -33.660 -158.600 ;
        RECT -32.460 -189.000 -0.600 -158.600 ;
        RECT 0.600 -189.000 32.460 -158.600 ;
        RECT 33.660 -189.000 65.520 -158.600 ;
        RECT 66.720 -189.000 98.580 -158.600 ;
        RECT 99.780 -189.000 131.640 -158.600 ;
        RECT 132.840 -189.000 164.700 -158.600 ;
        RECT 165.900 -189.000 197.760 -158.600 ;
      LAYER met4 ;
        RECT -182.820 188.605 -182.300 189.600 ;
        RECT -197.365 158.995 -167.755 188.605 ;
        RECT -182.820 157.005 -182.300 158.995 ;
        RECT -197.365 127.395 -167.755 157.005 ;
        RECT -182.820 125.405 -182.300 127.395 ;
        RECT -197.365 95.795 -167.755 125.405 ;
        RECT -182.820 93.805 -182.300 95.795 ;
        RECT -197.365 64.195 -167.755 93.805 ;
        RECT -182.820 62.205 -182.300 64.195 ;
        RECT -197.365 32.595 -167.755 62.205 ;
        RECT -182.820 30.605 -182.300 32.595 ;
        RECT -197.365 0.995 -167.755 30.605 ;
        RECT -182.820 -0.995 -182.300 0.995 ;
        RECT -197.365 -30.605 -167.755 -0.995 ;
        RECT -182.820 -32.595 -182.300 -30.605 ;
        RECT -197.365 -62.205 -167.755 -32.595 ;
        RECT -182.820 -64.195 -182.300 -62.205 ;
        RECT -197.365 -93.805 -167.755 -64.195 ;
        RECT -182.820 -95.795 -182.300 -93.805 ;
        RECT -197.365 -125.405 -167.755 -95.795 ;
        RECT -182.820 -127.395 -182.300 -125.405 ;
        RECT -197.365 -157.005 -167.755 -127.395 ;
        RECT -182.820 -158.995 -182.300 -157.005 ;
        RECT -197.365 -188.605 -167.755 -158.995 ;
        RECT -182.820 -189.600 -182.300 -188.605 ;
        RECT -166.420 -189.600 -165.900 189.600 ;
        RECT -149.760 188.605 -149.240 189.600 ;
        RECT -164.305 158.995 -134.695 188.605 ;
        RECT -149.760 157.005 -149.240 158.995 ;
        RECT -164.305 127.395 -134.695 157.005 ;
        RECT -149.760 125.405 -149.240 127.395 ;
        RECT -164.305 95.795 -134.695 125.405 ;
        RECT -149.760 93.805 -149.240 95.795 ;
        RECT -164.305 64.195 -134.695 93.805 ;
        RECT -149.760 62.205 -149.240 64.195 ;
        RECT -164.305 32.595 -134.695 62.205 ;
        RECT -149.760 30.605 -149.240 32.595 ;
        RECT -164.305 0.995 -134.695 30.605 ;
        RECT -149.760 -0.995 -149.240 0.995 ;
        RECT -164.305 -30.605 -134.695 -0.995 ;
        RECT -149.760 -32.595 -149.240 -30.605 ;
        RECT -164.305 -62.205 -134.695 -32.595 ;
        RECT -149.760 -64.195 -149.240 -62.205 ;
        RECT -164.305 -93.805 -134.695 -64.195 ;
        RECT -149.760 -95.795 -149.240 -93.805 ;
        RECT -164.305 -125.405 -134.695 -95.795 ;
        RECT -149.760 -127.395 -149.240 -125.405 ;
        RECT -164.305 -157.005 -134.695 -127.395 ;
        RECT -149.760 -158.995 -149.240 -157.005 ;
        RECT -164.305 -188.605 -134.695 -158.995 ;
        RECT -149.760 -189.600 -149.240 -188.605 ;
        RECT -133.360 -189.600 -132.840 189.600 ;
        RECT -116.700 188.605 -116.180 189.600 ;
        RECT -131.245 158.995 -101.635 188.605 ;
        RECT -116.700 157.005 -116.180 158.995 ;
        RECT -131.245 127.395 -101.635 157.005 ;
        RECT -116.700 125.405 -116.180 127.395 ;
        RECT -131.245 95.795 -101.635 125.405 ;
        RECT -116.700 93.805 -116.180 95.795 ;
        RECT -131.245 64.195 -101.635 93.805 ;
        RECT -116.700 62.205 -116.180 64.195 ;
        RECT -131.245 32.595 -101.635 62.205 ;
        RECT -116.700 30.605 -116.180 32.595 ;
        RECT -131.245 0.995 -101.635 30.605 ;
        RECT -116.700 -0.995 -116.180 0.995 ;
        RECT -131.245 -30.605 -101.635 -0.995 ;
        RECT -116.700 -32.595 -116.180 -30.605 ;
        RECT -131.245 -62.205 -101.635 -32.595 ;
        RECT -116.700 -64.195 -116.180 -62.205 ;
        RECT -131.245 -93.805 -101.635 -64.195 ;
        RECT -116.700 -95.795 -116.180 -93.805 ;
        RECT -131.245 -125.405 -101.635 -95.795 ;
        RECT -116.700 -127.395 -116.180 -125.405 ;
        RECT -131.245 -157.005 -101.635 -127.395 ;
        RECT -116.700 -158.995 -116.180 -157.005 ;
        RECT -131.245 -188.605 -101.635 -158.995 ;
        RECT -116.700 -189.600 -116.180 -188.605 ;
        RECT -100.300 -189.600 -99.780 189.600 ;
        RECT -83.640 188.605 -83.120 189.600 ;
        RECT -98.185 158.995 -68.575 188.605 ;
        RECT -83.640 157.005 -83.120 158.995 ;
        RECT -98.185 127.395 -68.575 157.005 ;
        RECT -83.640 125.405 -83.120 127.395 ;
        RECT -98.185 95.795 -68.575 125.405 ;
        RECT -83.640 93.805 -83.120 95.795 ;
        RECT -98.185 64.195 -68.575 93.805 ;
        RECT -83.640 62.205 -83.120 64.195 ;
        RECT -98.185 32.595 -68.575 62.205 ;
        RECT -83.640 30.605 -83.120 32.595 ;
        RECT -98.185 0.995 -68.575 30.605 ;
        RECT -83.640 -0.995 -83.120 0.995 ;
        RECT -98.185 -30.605 -68.575 -0.995 ;
        RECT -83.640 -32.595 -83.120 -30.605 ;
        RECT -98.185 -62.205 -68.575 -32.595 ;
        RECT -83.640 -64.195 -83.120 -62.205 ;
        RECT -98.185 -93.805 -68.575 -64.195 ;
        RECT -83.640 -95.795 -83.120 -93.805 ;
        RECT -98.185 -125.405 -68.575 -95.795 ;
        RECT -83.640 -127.395 -83.120 -125.405 ;
        RECT -98.185 -157.005 -68.575 -127.395 ;
        RECT -83.640 -158.995 -83.120 -157.005 ;
        RECT -98.185 -188.605 -68.575 -158.995 ;
        RECT -83.640 -189.600 -83.120 -188.605 ;
        RECT -67.240 -189.600 -66.720 189.600 ;
        RECT -50.580 188.605 -50.060 189.600 ;
        RECT -65.125 158.995 -35.515 188.605 ;
        RECT -50.580 157.005 -50.060 158.995 ;
        RECT -65.125 127.395 -35.515 157.005 ;
        RECT -50.580 125.405 -50.060 127.395 ;
        RECT -65.125 95.795 -35.515 125.405 ;
        RECT -50.580 93.805 -50.060 95.795 ;
        RECT -65.125 64.195 -35.515 93.805 ;
        RECT -50.580 62.205 -50.060 64.195 ;
        RECT -65.125 32.595 -35.515 62.205 ;
        RECT -50.580 30.605 -50.060 32.595 ;
        RECT -65.125 0.995 -35.515 30.605 ;
        RECT -50.580 -0.995 -50.060 0.995 ;
        RECT -65.125 -30.605 -35.515 -0.995 ;
        RECT -50.580 -32.595 -50.060 -30.605 ;
        RECT -65.125 -62.205 -35.515 -32.595 ;
        RECT -50.580 -64.195 -50.060 -62.205 ;
        RECT -65.125 -93.805 -35.515 -64.195 ;
        RECT -50.580 -95.795 -50.060 -93.805 ;
        RECT -65.125 -125.405 -35.515 -95.795 ;
        RECT -50.580 -127.395 -50.060 -125.405 ;
        RECT -65.125 -157.005 -35.515 -127.395 ;
        RECT -50.580 -158.995 -50.060 -157.005 ;
        RECT -65.125 -188.605 -35.515 -158.995 ;
        RECT -50.580 -189.600 -50.060 -188.605 ;
        RECT -34.180 -189.600 -33.660 189.600 ;
        RECT -17.520 188.605 -17.000 189.600 ;
        RECT -32.065 158.995 -2.455 188.605 ;
        RECT -17.520 157.005 -17.000 158.995 ;
        RECT -32.065 127.395 -2.455 157.005 ;
        RECT -17.520 125.405 -17.000 127.395 ;
        RECT -32.065 95.795 -2.455 125.405 ;
        RECT -17.520 93.805 -17.000 95.795 ;
        RECT -32.065 64.195 -2.455 93.805 ;
        RECT -17.520 62.205 -17.000 64.195 ;
        RECT -32.065 32.595 -2.455 62.205 ;
        RECT -17.520 30.605 -17.000 32.595 ;
        RECT -32.065 0.995 -2.455 30.605 ;
        RECT -17.520 -0.995 -17.000 0.995 ;
        RECT -32.065 -30.605 -2.455 -0.995 ;
        RECT -17.520 -32.595 -17.000 -30.605 ;
        RECT -32.065 -62.205 -2.455 -32.595 ;
        RECT -17.520 -64.195 -17.000 -62.205 ;
        RECT -32.065 -93.805 -2.455 -64.195 ;
        RECT -17.520 -95.795 -17.000 -93.805 ;
        RECT -32.065 -125.405 -2.455 -95.795 ;
        RECT -17.520 -127.395 -17.000 -125.405 ;
        RECT -32.065 -157.005 -2.455 -127.395 ;
        RECT -17.520 -158.995 -17.000 -157.005 ;
        RECT -32.065 -188.605 -2.455 -158.995 ;
        RECT -17.520 -189.600 -17.000 -188.605 ;
        RECT -1.120 -189.600 -0.600 189.600 ;
        RECT 15.540 188.605 16.060 189.600 ;
        RECT 0.995 158.995 30.605 188.605 ;
        RECT 15.540 157.005 16.060 158.995 ;
        RECT 0.995 127.395 30.605 157.005 ;
        RECT 15.540 125.405 16.060 127.395 ;
        RECT 0.995 95.795 30.605 125.405 ;
        RECT 15.540 93.805 16.060 95.795 ;
        RECT 0.995 64.195 30.605 93.805 ;
        RECT 15.540 62.205 16.060 64.195 ;
        RECT 0.995 32.595 30.605 62.205 ;
        RECT 15.540 30.605 16.060 32.595 ;
        RECT 0.995 0.995 30.605 30.605 ;
        RECT 15.540 -0.995 16.060 0.995 ;
        RECT 0.995 -30.605 30.605 -0.995 ;
        RECT 15.540 -32.595 16.060 -30.605 ;
        RECT 0.995 -62.205 30.605 -32.595 ;
        RECT 15.540 -64.195 16.060 -62.205 ;
        RECT 0.995 -93.805 30.605 -64.195 ;
        RECT 15.540 -95.795 16.060 -93.805 ;
        RECT 0.995 -125.405 30.605 -95.795 ;
        RECT 15.540 -127.395 16.060 -125.405 ;
        RECT 0.995 -157.005 30.605 -127.395 ;
        RECT 15.540 -158.995 16.060 -157.005 ;
        RECT 0.995 -188.605 30.605 -158.995 ;
        RECT 15.540 -189.600 16.060 -188.605 ;
        RECT 31.940 -189.600 32.460 189.600 ;
        RECT 48.600 188.605 49.120 189.600 ;
        RECT 34.055 158.995 63.665 188.605 ;
        RECT 48.600 157.005 49.120 158.995 ;
        RECT 34.055 127.395 63.665 157.005 ;
        RECT 48.600 125.405 49.120 127.395 ;
        RECT 34.055 95.795 63.665 125.405 ;
        RECT 48.600 93.805 49.120 95.795 ;
        RECT 34.055 64.195 63.665 93.805 ;
        RECT 48.600 62.205 49.120 64.195 ;
        RECT 34.055 32.595 63.665 62.205 ;
        RECT 48.600 30.605 49.120 32.595 ;
        RECT 34.055 0.995 63.665 30.605 ;
        RECT 48.600 -0.995 49.120 0.995 ;
        RECT 34.055 -30.605 63.665 -0.995 ;
        RECT 48.600 -32.595 49.120 -30.605 ;
        RECT 34.055 -62.205 63.665 -32.595 ;
        RECT 48.600 -64.195 49.120 -62.205 ;
        RECT 34.055 -93.805 63.665 -64.195 ;
        RECT 48.600 -95.795 49.120 -93.805 ;
        RECT 34.055 -125.405 63.665 -95.795 ;
        RECT 48.600 -127.395 49.120 -125.405 ;
        RECT 34.055 -157.005 63.665 -127.395 ;
        RECT 48.600 -158.995 49.120 -157.005 ;
        RECT 34.055 -188.605 63.665 -158.995 ;
        RECT 48.600 -189.600 49.120 -188.605 ;
        RECT 65.000 -189.600 65.520 189.600 ;
        RECT 81.660 188.605 82.180 189.600 ;
        RECT 67.115 158.995 96.725 188.605 ;
        RECT 81.660 157.005 82.180 158.995 ;
        RECT 67.115 127.395 96.725 157.005 ;
        RECT 81.660 125.405 82.180 127.395 ;
        RECT 67.115 95.795 96.725 125.405 ;
        RECT 81.660 93.805 82.180 95.795 ;
        RECT 67.115 64.195 96.725 93.805 ;
        RECT 81.660 62.205 82.180 64.195 ;
        RECT 67.115 32.595 96.725 62.205 ;
        RECT 81.660 30.605 82.180 32.595 ;
        RECT 67.115 0.995 96.725 30.605 ;
        RECT 81.660 -0.995 82.180 0.995 ;
        RECT 67.115 -30.605 96.725 -0.995 ;
        RECT 81.660 -32.595 82.180 -30.605 ;
        RECT 67.115 -62.205 96.725 -32.595 ;
        RECT 81.660 -64.195 82.180 -62.205 ;
        RECT 67.115 -93.805 96.725 -64.195 ;
        RECT 81.660 -95.795 82.180 -93.805 ;
        RECT 67.115 -125.405 96.725 -95.795 ;
        RECT 81.660 -127.395 82.180 -125.405 ;
        RECT 67.115 -157.005 96.725 -127.395 ;
        RECT 81.660 -158.995 82.180 -157.005 ;
        RECT 67.115 -188.605 96.725 -158.995 ;
        RECT 81.660 -189.600 82.180 -188.605 ;
        RECT 98.060 -189.600 98.580 189.600 ;
        RECT 114.720 188.605 115.240 189.600 ;
        RECT 100.175 158.995 129.785 188.605 ;
        RECT 114.720 157.005 115.240 158.995 ;
        RECT 100.175 127.395 129.785 157.005 ;
        RECT 114.720 125.405 115.240 127.395 ;
        RECT 100.175 95.795 129.785 125.405 ;
        RECT 114.720 93.805 115.240 95.795 ;
        RECT 100.175 64.195 129.785 93.805 ;
        RECT 114.720 62.205 115.240 64.195 ;
        RECT 100.175 32.595 129.785 62.205 ;
        RECT 114.720 30.605 115.240 32.595 ;
        RECT 100.175 0.995 129.785 30.605 ;
        RECT 114.720 -0.995 115.240 0.995 ;
        RECT 100.175 -30.605 129.785 -0.995 ;
        RECT 114.720 -32.595 115.240 -30.605 ;
        RECT 100.175 -62.205 129.785 -32.595 ;
        RECT 114.720 -64.195 115.240 -62.205 ;
        RECT 100.175 -93.805 129.785 -64.195 ;
        RECT 114.720 -95.795 115.240 -93.805 ;
        RECT 100.175 -125.405 129.785 -95.795 ;
        RECT 114.720 -127.395 115.240 -125.405 ;
        RECT 100.175 -157.005 129.785 -127.395 ;
        RECT 114.720 -158.995 115.240 -157.005 ;
        RECT 100.175 -188.605 129.785 -158.995 ;
        RECT 114.720 -189.600 115.240 -188.605 ;
        RECT 131.120 -189.600 131.640 189.600 ;
        RECT 147.780 188.605 148.300 189.600 ;
        RECT 133.235 158.995 162.845 188.605 ;
        RECT 147.780 157.005 148.300 158.995 ;
        RECT 133.235 127.395 162.845 157.005 ;
        RECT 147.780 125.405 148.300 127.395 ;
        RECT 133.235 95.795 162.845 125.405 ;
        RECT 147.780 93.805 148.300 95.795 ;
        RECT 133.235 64.195 162.845 93.805 ;
        RECT 147.780 62.205 148.300 64.195 ;
        RECT 133.235 32.595 162.845 62.205 ;
        RECT 147.780 30.605 148.300 32.595 ;
        RECT 133.235 0.995 162.845 30.605 ;
        RECT 147.780 -0.995 148.300 0.995 ;
        RECT 133.235 -30.605 162.845 -0.995 ;
        RECT 147.780 -32.595 148.300 -30.605 ;
        RECT 133.235 -62.205 162.845 -32.595 ;
        RECT 147.780 -64.195 148.300 -62.205 ;
        RECT 133.235 -93.805 162.845 -64.195 ;
        RECT 147.780 -95.795 148.300 -93.805 ;
        RECT 133.235 -125.405 162.845 -95.795 ;
        RECT 147.780 -127.395 148.300 -125.405 ;
        RECT 133.235 -157.005 162.845 -127.395 ;
        RECT 147.780 -158.995 148.300 -157.005 ;
        RECT 133.235 -188.605 162.845 -158.995 ;
        RECT 147.780 -189.600 148.300 -188.605 ;
        RECT 164.180 -189.600 164.700 189.600 ;
        RECT 180.840 188.605 181.360 189.600 ;
        RECT 166.295 158.995 195.905 188.605 ;
        RECT 180.840 157.005 181.360 158.995 ;
        RECT 166.295 127.395 195.905 157.005 ;
        RECT 180.840 125.405 181.360 127.395 ;
        RECT 166.295 95.795 195.905 125.405 ;
        RECT 180.840 93.805 181.360 95.795 ;
        RECT 166.295 64.195 195.905 93.805 ;
        RECT 180.840 62.205 181.360 64.195 ;
        RECT 166.295 32.595 195.905 62.205 ;
        RECT 180.840 30.605 181.360 32.595 ;
        RECT 166.295 0.995 195.905 30.605 ;
        RECT 180.840 -0.995 181.360 0.995 ;
        RECT 166.295 -30.605 195.905 -0.995 ;
        RECT 180.840 -32.595 181.360 -30.605 ;
        RECT 166.295 -62.205 195.905 -32.595 ;
        RECT 180.840 -64.195 181.360 -62.205 ;
        RECT 166.295 -93.805 195.905 -64.195 ;
        RECT 180.840 -95.795 181.360 -93.805 ;
        RECT 166.295 -125.405 195.905 -95.795 ;
        RECT 180.840 -127.395 181.360 -125.405 ;
        RECT 166.295 -157.005 195.905 -127.395 ;
        RECT 180.840 -158.995 181.360 -157.005 ;
        RECT 166.295 -188.605 195.905 -158.995 ;
        RECT 180.840 -189.600 181.360 -188.605 ;
        RECT 197.240 -189.600 197.760 189.600 ;
  END
END sky130_fd_pr__cap_mim_m3_1_Z926RQ
MACRO sky130_fd_pr__cap_mim_m3_1_39XMLG
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__cap_mim_m3_1_39XMLG ;
  ORIGIN -50.190 -48.000 ;
  SIZE 30.400 BY 30.400 ;
  OBS
      LAYER met3 ;
        RECT -82.050 48.000 -50.190 78.400 ;
        RECT -48.990 48.000 -17.130 78.400 ;
        RECT -15.930 48.000 15.930 78.400 ;
        RECT 17.130 48.000 48.990 78.400 ;
        RECT 50.190 48.000 82.050 78.400 ;
        RECT -82.050 16.400 -50.190 46.800 ;
        RECT -48.990 16.400 -17.130 46.800 ;
        RECT -15.930 16.400 15.930 46.800 ;
        RECT 17.130 16.400 48.990 46.800 ;
        RECT 50.190 16.400 82.050 46.800 ;
        RECT -82.050 -15.200 -50.190 15.200 ;
        RECT -48.990 -15.200 -17.130 15.200 ;
        RECT -15.930 -15.200 15.930 15.200 ;
        RECT 17.130 -15.200 48.990 15.200 ;
        RECT 50.190 -15.200 82.050 15.200 ;
        RECT -82.050 -46.800 -50.190 -16.400 ;
        RECT -48.990 -46.800 -17.130 -16.400 ;
        RECT -15.930 -46.800 15.930 -16.400 ;
        RECT 17.130 -46.800 48.990 -16.400 ;
        RECT 50.190 -46.800 82.050 -16.400 ;
        RECT -82.050 -78.400 -50.190 -48.000 ;
        RECT -48.990 -78.400 -17.130 -48.000 ;
        RECT -15.930 -78.400 15.930 -48.000 ;
        RECT 17.130 -78.400 48.990 -48.000 ;
        RECT 50.190 -78.400 82.050 -48.000 ;
      LAYER met4 ;
        RECT -67.110 78.005 -66.590 79.000 ;
        RECT -81.655 48.395 -52.045 78.005 ;
        RECT -67.110 46.405 -66.590 48.395 ;
        RECT -81.655 16.795 -52.045 46.405 ;
        RECT -67.110 14.805 -66.590 16.795 ;
        RECT -81.655 -14.805 -52.045 14.805 ;
        RECT -67.110 -16.795 -66.590 -14.805 ;
        RECT -81.655 -46.405 -52.045 -16.795 ;
        RECT -67.110 -48.395 -66.590 -46.405 ;
        RECT -81.655 -78.005 -52.045 -48.395 ;
        RECT -67.110 -79.000 -66.590 -78.005 ;
        RECT -50.710 -79.000 -50.190 79.000 ;
        RECT -34.050 78.005 -33.530 79.000 ;
        RECT -48.595 48.395 -18.985 78.005 ;
        RECT -34.050 46.405 -33.530 48.395 ;
        RECT -48.595 16.795 -18.985 46.405 ;
        RECT -34.050 14.805 -33.530 16.795 ;
        RECT -48.595 -14.805 -18.985 14.805 ;
        RECT -34.050 -16.795 -33.530 -14.805 ;
        RECT -48.595 -46.405 -18.985 -16.795 ;
        RECT -34.050 -48.395 -33.530 -46.405 ;
        RECT -48.595 -78.005 -18.985 -48.395 ;
        RECT -34.050 -79.000 -33.530 -78.005 ;
        RECT -17.650 -79.000 -17.130 79.000 ;
        RECT -0.990 78.005 -0.470 79.000 ;
        RECT -15.535 48.395 14.075 78.005 ;
        RECT -0.990 46.405 -0.470 48.395 ;
        RECT -15.535 16.795 14.075 46.405 ;
        RECT -0.990 14.805 -0.470 16.795 ;
        RECT -15.535 -14.805 14.075 14.805 ;
        RECT -0.990 -16.795 -0.470 -14.805 ;
        RECT -15.535 -46.405 14.075 -16.795 ;
        RECT -0.990 -48.395 -0.470 -46.405 ;
        RECT -15.535 -78.005 14.075 -48.395 ;
        RECT -0.990 -79.000 -0.470 -78.005 ;
        RECT 15.410 -79.000 15.930 79.000 ;
        RECT 32.070 78.005 32.590 79.000 ;
        RECT 17.525 48.395 47.135 78.005 ;
        RECT 32.070 46.405 32.590 48.395 ;
        RECT 17.525 16.795 47.135 46.405 ;
        RECT 32.070 14.805 32.590 16.795 ;
        RECT 17.525 -14.805 47.135 14.805 ;
        RECT 32.070 -16.795 32.590 -14.805 ;
        RECT 17.525 -46.405 47.135 -16.795 ;
        RECT 32.070 -48.395 32.590 -46.405 ;
        RECT 17.525 -78.005 47.135 -48.395 ;
        RECT 32.070 -79.000 32.590 -78.005 ;
        RECT 48.470 -79.000 48.990 79.000 ;
        RECT 65.130 78.005 65.650 79.000 ;
        RECT 50.585 48.395 80.195 78.005 ;
        RECT 65.130 46.405 65.650 48.395 ;
        RECT 50.585 16.795 80.195 46.405 ;
        RECT 65.130 14.805 65.650 16.795 ;
        RECT 50.585 -14.805 80.195 14.805 ;
        RECT 65.130 -16.795 65.650 -14.805 ;
        RECT 50.585 -46.405 80.195 -16.795 ;
        RECT 65.130 -48.395 65.650 -46.405 ;
        RECT 50.585 -78.005 80.195 -48.395 ;
        RECT 65.130 -79.000 65.650 -78.005 ;
        RECT 81.530 -79.000 82.050 79.000 ;
  END
END sky130_fd_pr__cap_mim_m3_1_39XMLG
MACRO sky130_fd_pr__res_generic_po_447X6E
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__res_generic_po_447X6E ;
  ORIGIN 0.805 3.540 ;
  SIZE 1.610 BY 7.080 ;
  OBS
      LAYER pwell ;
        RECT -1.070 -3.805 1.070 3.805 ;
      LAYER li1 ;
        RECT -0.890 3.455 0.890 3.625 ;
        RECT -0.890 -3.455 -0.720 3.455 ;
        RECT -0.240 2.725 0.240 2.895 ;
        RECT -0.160 0.910 0.160 2.725 ;
        RECT -0.160 -2.725 0.160 -0.910 ;
        RECT -0.240 -2.895 0.240 -2.725 ;
        RECT 0.720 -3.455 0.890 3.455 ;
        RECT -0.890 -3.625 0.890 -3.455 ;
      LAYER met1 ;
        RECT -0.190 0.850 0.190 2.955 ;
        RECT -0.190 -2.955 0.190 -0.850 ;
  END
END sky130_fd_pr__res_generic_po_447X6E
MACRO sky130_fd_pr__pfet_01v8_7PMXFU
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_7PMXFU ;
  ORIGIN 0.805 23.330 ;
  SIZE 1.610 BY 46.660 ;
  OBS
      LAYER nwell ;
        RECT -1.070 -23.595 1.070 23.595 ;
      LAYER li1 ;
        RECT -0.890 23.245 0.890 23.415 ;
        RECT -0.890 -23.245 -0.720 23.245 ;
        RECT -0.165 22.735 0.165 22.905 ;
        RECT -0.320 -22.520 -0.150 22.520 ;
        RECT 0.150 -22.520 0.320 22.520 ;
        RECT -0.165 -22.905 0.165 -22.735 ;
        RECT 0.720 -23.245 0.890 23.245 ;
        RECT -0.890 -23.415 0.890 -23.245 ;
      LAYER met1 ;
        RECT -0.780 23.215 0.780 23.445 ;
        RECT -0.145 22.705 0.145 22.935 ;
        RECT -0.350 4.345 -0.120 22.415 ;
        RECT 0.120 -22.415 0.350 -4.345 ;
        RECT -0.145 -22.935 0.145 -22.705 ;
  END
END sky130_fd_pr__pfet_01v8_7PMXFU
MACRO sky130_fd_pr__pfet_01v8_KXJ7FM
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_KXJ7FM ;
  ORIGIN 0.805 1.100 ;
  SIZE 1.610 BY 2.200 ;
  OBS
      LAYER nwell ;
        RECT -1.070 -1.365 1.070 1.365 ;
      LAYER li1 ;
        RECT -0.890 1.015 0.890 1.185 ;
        RECT -0.890 -1.015 -0.720 1.015 ;
        RECT -0.165 0.505 0.165 0.675 ;
        RECT -0.320 -0.290 -0.150 0.290 ;
        RECT 0.150 -0.290 0.320 0.290 ;
        RECT -0.165 -0.675 0.165 -0.505 ;
        RECT 0.720 -1.015 0.890 1.015 ;
        RECT -0.890 -1.185 0.890 -1.015 ;
      LAYER met1 ;
        RECT 0.085 0.985 0.780 1.215 ;
        RECT -0.145 0.475 0.145 0.705 ;
        RECT -0.350 -0.270 -0.120 0.270 ;
        RECT 0.120 -0.270 0.350 0.270 ;
        RECT -0.145 -0.705 0.145 -0.475 ;
  END
END sky130_fd_pr__pfet_01v8_KXJ7FM
MACRO sky130_fd_pr__pfet_01v8_K9S5FM
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_K9S5FM ;
  ORIGIN 0.805 1.100 ;
  SIZE 1.610 BY 2.200 ;
  OBS
      LAYER nwell ;
        RECT -1.070 -1.365 1.070 1.365 ;
      LAYER li1 ;
        RECT -0.890 1.015 0.890 1.185 ;
        RECT -0.890 -1.015 -0.720 1.015 ;
        RECT -0.165 0.505 0.165 0.675 ;
        RECT -0.320 -0.290 -0.150 0.290 ;
        RECT 0.150 -0.290 0.320 0.290 ;
        RECT -0.165 -0.675 0.165 -0.505 ;
        RECT 0.720 -1.015 0.890 1.015 ;
        RECT -0.890 -1.185 0.890 -1.015 ;
      LAYER met1 ;
        RECT -0.145 0.475 0.145 0.705 ;
        RECT -0.350 -0.270 -0.120 0.270 ;
        RECT 0.120 -0.270 0.350 0.270 ;
        RECT -0.145 -0.705 0.145 -0.475 ;
        RECT 0.690 -1.075 0.920 1.075 ;
  END
END sky130_fd_pr__pfet_01v8_K9S5FM
MACRO sky130_fd_pr__pfet_01v8_K9S7EM
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_K9S7EM ;
  ORIGIN 0.805 1.100 ;
  SIZE 1.610 BY 2.200 ;
  OBS
      LAYER nwell ;
        RECT -1.070 -1.365 1.070 1.365 ;
      LAYER li1 ;
        RECT -0.890 1.015 0.890 1.185 ;
        RECT -0.890 -1.015 -0.720 1.015 ;
        RECT -0.165 0.505 0.165 0.675 ;
        RECT -0.320 -0.290 -0.150 0.290 ;
        RECT 0.150 -0.290 0.320 0.290 ;
        RECT -0.165 -0.675 0.165 -0.505 ;
        RECT 0.720 -1.015 0.890 1.015 ;
        RECT -0.890 -1.185 0.890 -1.015 ;
      LAYER met1 ;
        RECT -0.145 0.475 0.145 0.705 ;
        RECT -0.350 -0.270 -0.120 0.270 ;
        RECT 0.120 -0.270 0.350 0.270 ;
        RECT -0.145 -0.705 0.145 -0.475 ;
        RECT -0.780 -1.215 0.780 -0.985 ;
  END
END sky130_fd_pr__pfet_01v8_K9S7EM
MACRO sky130_fd_pr__pfet_01v8_KZR7FM
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_KZR7FM ;
  ORIGIN 0.805 1.100 ;
  SIZE 1.610 BY 2.200 ;
  OBS
      LAYER nwell ;
        RECT -1.070 -1.365 1.070 1.365 ;
      LAYER li1 ;
        RECT -0.890 1.015 0.890 1.185 ;
        RECT -0.890 -1.015 -0.720 1.015 ;
        RECT -0.165 0.505 0.165 0.675 ;
        RECT -0.320 -0.290 -0.150 0.290 ;
        RECT 0.150 -0.290 0.320 0.290 ;
        RECT -0.165 -0.675 0.165 -0.505 ;
        RECT 0.720 -1.015 0.890 1.015 ;
        RECT -0.890 -1.185 0.890 -1.015 ;
      LAYER met1 ;
        RECT -0.780 0.985 0.780 1.215 ;
        RECT -0.145 0.475 0.145 0.705 ;
        RECT -0.350 -0.270 -0.120 0.270 ;
        RECT 0.120 -0.270 0.350 0.270 ;
        RECT -0.145 -0.705 0.145 -0.475 ;
  END
END sky130_fd_pr__pfet_01v8_KZR7FM
MACRO sky130_fd_pr__nfet_01v8_6FB27G
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__nfet_01v8_6FB27G ;
  ORIGIN 0.805 0.995 ;
  SIZE 1.610 BY 1.990 ;
  OBS
      LAYER pwell ;
        RECT -1.070 -1.260 1.070 1.260 ;
      LAYER li1 ;
        RECT -0.890 0.910 0.890 1.080 ;
        RECT -0.890 -0.910 -0.720 0.910 ;
        RECT -0.165 0.400 0.165 0.570 ;
        RECT -0.320 -0.230 -0.150 0.230 ;
        RECT 0.150 -0.230 0.320 0.230 ;
        RECT -0.165 -0.570 0.165 -0.400 ;
        RECT 0.720 -0.910 0.890 0.910 ;
        RECT -0.890 -1.080 0.890 -0.910 ;
      LAYER met1 ;
        RECT -0.145 0.370 0.145 0.600 ;
        RECT -0.350 -0.210 -0.120 0.210 ;
        RECT 0.120 -0.210 0.350 0.210 ;
        RECT -0.145 -0.600 0.145 -0.370 ;
        RECT 0.690 -0.970 0.920 0.970 ;
  END
END sky130_fd_pr__nfet_01v8_6FB27G
MACRO sky130_fd_pr__nfet_01v8_6FB46G
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__nfet_01v8_6FB46G ;
  ORIGIN 0.805 0.995 ;
  SIZE 1.610 BY 1.990 ;
  OBS
      LAYER pwell ;
        RECT -1.070 -1.260 1.070 1.260 ;
      LAYER li1 ;
        RECT -0.890 0.910 0.890 1.080 ;
        RECT -0.890 -0.910 -0.720 0.910 ;
        RECT -0.165 0.400 0.165 0.570 ;
        RECT -0.320 -0.230 -0.150 0.230 ;
        RECT 0.150 -0.230 0.320 0.230 ;
        RECT -0.165 -0.570 0.165 -0.400 ;
        RECT 0.720 -0.910 0.890 0.910 ;
        RECT -0.890 -1.080 0.890 -0.910 ;
      LAYER met1 ;
        RECT -0.145 0.370 0.145 0.600 ;
        RECT -0.350 -0.210 -0.120 0.210 ;
        RECT 0.120 -0.210 0.350 0.210 ;
        RECT -0.145 -0.600 0.145 -0.370 ;
        RECT -0.780 -1.110 0.780 -0.880 ;
  END
END sky130_fd_pr__nfet_01v8_6FB46G
MACRO sky130_fd_pr__nfet_01v8_HAAXKC
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__nfet_01v8_HAAXKC ;
  ORIGIN 0.805 8.285 ;
  SIZE 1.610 BY 16.570 ;
  OBS
      LAYER pwell ;
        RECT -1.070 -8.550 1.070 8.550 ;
      LAYER li1 ;
        RECT -0.890 8.200 0.890 8.370 ;
        RECT -0.890 -8.200 -0.720 8.200 ;
        RECT -0.165 7.690 0.165 7.860 ;
        RECT -0.320 -7.520 -0.150 7.520 ;
        RECT 0.150 -7.520 0.320 7.520 ;
        RECT -0.165 -7.860 0.165 -7.690 ;
        RECT 0.720 -8.200 0.890 8.200 ;
        RECT -0.890 -8.370 0.890 -8.200 ;
      LAYER met1 ;
        RECT -0.145 7.660 0.145 7.890 ;
        RECT -0.350 1.345 -0.120 7.415 ;
        RECT 0.120 -7.415 0.350 -1.345 ;
        RECT -0.145 -7.890 0.145 -7.660 ;
        RECT -0.780 -8.400 0.780 -8.170 ;
  END
END sky130_fd_pr__nfet_01v8_HAAXKC
MACRO cp
  CLASS BLOCK ;
  FOREIGN cp ;
  ORIGIN 327.630 5.190 ;
  SIZE 586.465 BY 447.700 ;
  PIN up
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.185 27.370 2.515 27.540 ;
        RECT 2.185 26.190 2.515 26.360 ;
        RECT 2.205 24.430 2.535 24.600 ;
        RECT 2.205 23.460 2.535 23.630 ;
        RECT 18.445 19.800 18.775 19.970 ;
        RECT 18.445 18.620 18.775 18.790 ;
      LAYER met1 ;
        RECT -0.380 27.350 2.530 27.580 ;
        RECT -0.380 26.375 -0.150 27.350 ;
        RECT 2.205 27.340 2.495 27.350 ;
        RECT 2.205 26.375 2.495 26.390 ;
        RECT -0.380 26.160 2.495 26.375 ;
        RECT -0.380 26.145 2.485 26.160 ;
        RECT -2.430 25.490 -1.430 25.860 ;
        RECT -0.380 25.490 -0.150 26.145 ;
        RECT -2.430 25.270 -0.150 25.490 ;
        RECT -2.430 24.860 -1.430 25.270 ;
        RECT -0.940 18.200 -0.720 25.270 ;
        RECT -0.380 24.665 -0.150 25.270 ;
        RECT -0.380 24.435 2.525 24.665 ;
        RECT -0.380 23.645 -0.150 24.435 ;
        RECT 2.225 24.400 2.515 24.435 ;
        RECT 2.225 23.645 2.515 23.660 ;
        RECT -0.380 23.415 2.525 23.645 ;
        RECT 16.020 20.000 18.740 20.010 ;
        RECT 16.020 19.790 18.755 20.000 ;
        RECT 16.020 18.770 16.240 19.790 ;
        RECT 18.465 19.770 18.755 19.790 ;
        RECT 18.465 18.770 18.755 18.820 ;
        RECT 16.000 18.550 18.780 18.770 ;
        RECT 1.540 18.200 1.860 18.220 ;
        RECT -0.940 17.980 1.860 18.200 ;
        RECT 1.540 17.960 1.860 17.980 ;
        RECT 3.070 18.200 3.330 18.250 ;
        RECT 5.880 18.200 6.200 18.220 ;
        RECT 3.070 17.980 6.200 18.200 ;
        RECT 3.070 17.930 3.330 17.980 ;
        RECT 5.880 17.960 6.200 17.980 ;
        RECT 7.730 18.200 7.990 18.250 ;
        RECT 16.000 18.200 16.220 18.550 ;
        RECT 7.730 17.980 16.220 18.200 ;
        RECT 7.730 17.930 7.990 17.980 ;
      LAYER met2 ;
        RECT 1.570 18.200 1.830 18.250 ;
        RECT 3.040 18.200 3.360 18.220 ;
        RECT 1.570 17.980 3.360 18.200 ;
        RECT 1.570 17.930 1.830 17.980 ;
        RECT 3.040 17.960 3.360 17.980 ;
        RECT 5.910 18.200 6.170 18.250 ;
        RECT 7.700 18.200 8.020 18.220 ;
        RECT 5.910 17.980 8.020 18.200 ;
        RECT 5.910 17.930 6.170 17.980 ;
        RECT 7.700 17.960 8.020 17.980 ;
    END
  END up
  PIN vctrl
    ANTENNADIFFAREA 0.278400 ;
    PORT
      LAYER li1 ;
        RECT 57.600 37.150 57.920 38.965 ;
        RECT 57.520 36.980 58.000 37.150 ;
        RECT 26.650 26.495 26.820 27.075 ;
        RECT 33.920 12.680 34.090 13.140 ;
      LAYER met1 ;
        RECT 74.680 98.020 85.450 98.460 ;
        RECT 57.570 36.920 57.950 39.025 ;
        RECT 57.600 35.870 57.920 36.920 ;
        RECT 57.600 35.520 57.900 35.870 ;
        RECT 57.560 35.080 57.900 35.520 ;
        RECT 57.600 34.680 57.900 35.080 ;
        RECT 57.600 29.720 57.920 34.680 ;
        RECT 36.710 29.400 57.920 29.720 ;
        RECT 26.620 26.920 26.850 27.055 ;
        RECT 26.620 26.710 28.210 26.920 ;
        RECT 26.620 26.515 26.850 26.710 ;
        RECT 28.000 21.020 28.210 26.710 ;
        RECT 36.710 21.020 37.030 29.400 ;
        RECT 74.680 24.120 75.120 98.020 ;
        RECT 40.530 23.680 75.120 24.120 ;
        RECT 40.530 21.020 40.970 23.680 ;
        RECT 44.960 21.020 45.960 21.530 ;
        RECT 27.970 20.660 45.960 21.020 ;
        RECT 28.000 14.295 28.210 20.660 ;
        RECT 44.960 20.210 45.960 20.660 ;
        RECT 32.790 14.295 33.110 14.320 ;
        RECT 28.000 14.085 33.110 14.295 ;
        RECT 32.790 14.060 33.110 14.085 ;
        RECT 32.790 13.005 33.110 13.030 ;
        RECT 33.890 13.005 34.120 13.120 ;
        RECT 32.790 12.795 34.120 13.005 ;
        RECT 32.790 12.770 33.110 12.795 ;
        RECT 33.890 12.700 34.120 12.795 ;
      LAYER met2 ;
        RECT 84.980 98.460 85.420 98.490 ;
        RECT 84.980 98.020 87.095 98.460 ;
        RECT 84.980 97.990 85.420 98.020 ;
        RECT 32.820 14.030 33.080 14.350 ;
        RECT 32.845 13.060 33.055 14.030 ;
        RECT 32.820 12.740 33.080 13.060 ;
      LAYER met3 ;
        RECT 255.990 183.000 256.570 183.520 ;
        RECT 256.020 179.195 256.540 183.000 ;
        RECT 255.995 178.685 256.565 179.195 ;
        RECT 256.020 178.680 256.540 178.685 ;
        RECT 86.585 98.460 87.075 98.485 ;
        RECT 86.585 98.020 88.890 98.460 ;
        RECT 86.585 97.995 87.075 98.020 ;
      LAYER met4 ;
        RECT 98.225 230.720 127.835 245.265 ;
        RECT 129.825 230.720 159.435 245.265 ;
        RECT 161.425 230.720 191.035 245.265 ;
        RECT 193.025 230.720 222.635 245.265 ;
        RECT 224.625 230.720 254.235 245.265 ;
        RECT 97.230 230.710 255.230 230.720 ;
        RECT 95.100 230.200 255.230 230.710 ;
        RECT 95.100 230.190 127.835 230.200 ;
        RECT 95.100 197.660 95.620 230.190 ;
        RECT 98.225 215.655 127.835 230.190 ;
        RECT 129.825 215.655 159.435 230.200 ;
        RECT 161.425 215.655 191.035 230.200 ;
        RECT 193.025 215.655 222.635 230.200 ;
        RECT 224.625 215.655 254.235 230.200 ;
        RECT 98.225 197.660 127.835 212.205 ;
        RECT 129.825 197.660 159.435 212.205 ;
        RECT 161.425 197.660 191.035 212.205 ;
        RECT 193.025 197.660 222.635 212.205 ;
        RECT 224.625 197.660 254.235 212.205 ;
        RECT 254.820 197.660 256.540 197.680 ;
        RECT 95.100 197.160 256.540 197.660 ;
        RECT 95.100 197.140 255.230 197.160 ;
        RECT 98.225 182.595 127.835 197.140 ;
        RECT 129.825 182.595 159.435 197.140 ;
        RECT 161.425 182.595 191.035 197.140 ;
        RECT 193.025 182.595 222.635 197.140 ;
        RECT 224.625 182.595 254.235 197.140 ;
        RECT 256.020 183.525 256.540 197.160 ;
        RECT 256.015 182.995 256.545 183.525 ;
        RECT 98.225 164.600 127.835 179.145 ;
        RECT 129.825 164.600 159.435 179.145 ;
        RECT 161.425 164.600 191.035 179.145 ;
        RECT 193.025 164.600 222.635 179.145 ;
        RECT 224.625 164.600 254.235 179.145 ;
        RECT 256.020 164.600 256.540 179.200 ;
        RECT 97.230 164.590 256.540 164.600 ;
        RECT 93.500 164.080 256.540 164.590 ;
        RECT 93.500 164.070 97.770 164.080 ;
        RECT 93.500 131.540 94.020 164.070 ;
        RECT 98.225 149.535 127.835 164.080 ;
        RECT 129.825 149.535 159.435 164.080 ;
        RECT 161.425 149.535 191.035 164.080 ;
        RECT 193.025 149.535 222.635 164.080 ;
        RECT 224.625 149.535 254.235 164.080 ;
        RECT 98.225 131.540 127.835 146.085 ;
        RECT 129.825 131.540 159.435 146.085 ;
        RECT 161.425 131.540 191.035 146.085 ;
        RECT 193.025 131.540 222.635 146.085 ;
        RECT 224.625 131.540 254.235 146.085 ;
        RECT 255.040 131.540 257.080 131.600 ;
        RECT 93.500 131.080 257.080 131.540 ;
        RECT 93.500 131.020 255.230 131.080 ;
        RECT 98.225 116.475 127.835 131.020 ;
        RECT 129.825 116.475 159.435 131.020 ;
        RECT 161.425 116.475 191.035 131.020 ;
        RECT 193.025 116.475 222.635 131.020 ;
        RECT 224.625 116.475 254.235 131.020 ;
        RECT 98.225 98.480 127.835 113.025 ;
        RECT 129.825 98.480 159.435 113.025 ;
        RECT 161.425 98.480 191.035 113.025 ;
        RECT 193.025 98.480 222.635 113.025 ;
        RECT 224.625 98.480 254.235 113.025 ;
        RECT 256.560 98.480 257.080 131.080 ;
        RECT 88.415 98.460 88.865 98.465 ;
        RECT 97.230 98.460 257.080 98.480 ;
        RECT 88.415 98.020 257.080 98.460 ;
        RECT 88.415 98.015 88.865 98.020 ;
        RECT 97.230 97.960 257.080 98.020 ;
        RECT 98.225 83.415 127.835 97.960 ;
        RECT 129.825 83.415 159.435 97.960 ;
        RECT 161.425 83.415 191.035 97.960 ;
        RECT 193.025 83.415 222.635 97.960 ;
        RECT 224.625 83.415 254.235 97.960 ;
    END
  END vctrl
  PIN VDD
    ANTENNAGATEAREA 0.345600 ;
    ANTENNADIFFAREA 33.939598 ;
    PORT
      LAYER nwell ;
        RECT -5.790 32.030 41.400 34.170 ;
        RECT 1.280 25.500 3.420 28.230 ;
        RECT 19.720 25.300 21.860 28.030 ;
        RECT 1.940 11.700 4.080 14.430 ;
      LAYER li1 ;
        RECT -5.610 33.820 41.220 33.990 ;
        RECT -5.610 32.380 -5.440 33.820 ;
        RECT -4.715 33.250 40.325 33.420 ;
        RECT 41.050 32.380 41.220 33.820 ;
        RECT -5.610 32.210 41.220 32.380 ;
        RECT 1.460 27.880 3.240 28.050 ;
        RECT 1.460 25.850 1.630 27.880 ;
        RECT 2.030 26.575 2.200 27.155 ;
        RECT 3.070 25.850 3.240 27.880 ;
        RECT 19.900 27.680 21.680 27.850 ;
        RECT 10.315 27.420 10.645 27.590 ;
        RECT 10.315 26.240 10.645 26.410 ;
        RECT 1.460 25.680 3.240 25.850 ;
        RECT 19.900 25.650 20.070 27.680 ;
        RECT 20.940 26.375 21.110 26.955 ;
        RECT 21.510 25.650 21.680 27.680 ;
        RECT 19.900 25.480 21.680 25.650 ;
        RECT 2.120 14.080 3.900 14.250 ;
        RECT 23.675 14.090 24.005 14.260 ;
        RECT 2.120 12.050 2.290 14.080 ;
        RECT 2.690 12.775 2.860 13.355 ;
        RECT 3.730 12.050 3.900 14.080 ;
        RECT 11.205 13.640 11.535 13.810 ;
        RECT 23.990 13.460 24.160 13.920 ;
        RECT 34.075 13.310 34.405 13.480 ;
        RECT 23.675 13.120 24.005 13.290 ;
        RECT 11.205 12.460 11.535 12.630 ;
        RECT 34.075 12.340 34.405 12.510 ;
        RECT 2.120 11.880 3.900 12.050 ;
      LAYER met1 ;
        RECT 39.120 34.745 39.350 34.790 ;
        RECT 39.120 34.515 41.795 34.745 ;
        RECT 39.120 33.450 39.350 34.515 ;
        RECT 41.565 34.050 41.795 34.515 ;
        RECT 22.150 33.220 40.220 33.450 ;
        RECT 40.980 32.230 41.990 34.050 ;
        RECT 41.425 30.905 41.755 32.230 ;
        RECT 33.755 30.575 41.755 30.905 ;
        RECT 19.220 30.195 19.550 30.210 ;
        RECT 26.535 30.195 26.865 30.225 ;
        RECT 33.755 30.195 34.085 30.575 ;
        RECT 8.850 29.720 9.850 30.110 ;
        RECT -3.750 29.370 9.850 29.720 ;
        RECT -3.750 15.365 -3.400 29.370 ;
        RECT 8.850 29.000 9.850 29.370 ;
        RECT 19.220 29.865 22.815 30.195 ;
        RECT 26.535 29.865 34.085 30.195 ;
        RECT 19.220 29.260 19.550 29.865 ;
        RECT 26.535 29.835 26.865 29.865 ;
        RECT 19.050 29.000 19.550 29.260 ;
        RECT 1.400 28.970 19.550 29.000 ;
        RECT 1.400 28.450 19.630 28.970 ;
        RECT 0.640 28.070 0.960 28.100 ;
        RECT 1.490 28.070 3.350 28.450 ;
        RECT 0.640 27.880 3.350 28.070 ;
        RECT 0.640 27.870 3.130 27.880 ;
        RECT 0.640 27.840 0.960 27.870 ;
        RECT 1.570 27.850 3.130 27.870 ;
        RECT 8.320 27.620 8.600 28.450 ;
        RECT 19.235 28.345 19.630 28.450 ;
        RECT 21.660 28.345 21.980 28.370 ;
        RECT 19.235 28.135 21.980 28.345 ;
        RECT 20.195 27.880 20.405 28.135 ;
        RECT 21.660 28.110 21.980 28.135 ;
        RECT 20.010 27.650 21.570 27.880 ;
        RECT 8.300 27.360 10.640 27.620 ;
        RECT 8.300 27.260 8.600 27.360 ;
        RECT 0.640 26.990 0.960 27.020 ;
        RECT 2.000 26.990 2.230 27.135 ;
        RECT 0.640 26.790 2.230 26.990 ;
        RECT 0.640 26.760 0.960 26.790 ;
        RECT 2.000 26.595 2.230 26.790 ;
        RECT 8.300 26.160 8.560 27.260 ;
        RECT 20.910 26.770 21.140 26.935 ;
        RECT 21.660 26.770 21.980 26.795 ;
        RECT 20.910 26.560 21.980 26.770 ;
        RECT 9.490 26.450 9.750 26.480 ;
        RECT 9.490 26.190 10.650 26.450 ;
        RECT 20.910 26.395 21.140 26.560 ;
        RECT 21.660 26.535 21.980 26.560 ;
        RECT 9.490 26.160 9.750 26.190 ;
        RECT -0.725 15.885 -0.375 15.915 ;
        RECT 7.020 15.885 8.020 16.020 ;
        RECT -0.725 15.535 8.020 15.885 ;
        RECT -0.725 15.505 -0.375 15.535 ;
        RECT -3.780 15.015 -3.370 15.365 ;
        RECT 7.020 15.010 8.020 15.535 ;
        RECT 16.095 15.105 26.535 15.335 ;
        RECT 2.360 14.860 15.220 15.010 ;
        RECT 2.240 14.855 15.220 14.860 ;
        RECT 16.095 14.855 16.325 15.105 ;
        RECT 2.240 14.840 16.325 14.855 ;
        RECT 1.740 14.640 16.325 14.840 ;
        RECT 1.740 14.270 1.940 14.640 ;
        RECT 2.240 14.625 16.325 14.640 ;
        RECT 2.240 14.580 15.220 14.625 ;
        RECT 2.240 14.280 4.120 14.580 ;
        RECT 1.680 14.010 2.000 14.270 ;
        RECT 2.230 14.110 4.120 14.280 ;
        RECT 2.230 14.050 3.790 14.110 ;
        RECT 8.390 13.680 8.670 14.580 ;
        RECT 26.305 14.395 26.535 15.105 ;
        RECT 23.735 14.290 26.945 14.395 ;
        RECT 23.695 14.165 26.945 14.290 ;
        RECT 23.695 14.060 23.985 14.165 ;
        RECT 23.960 13.840 24.190 13.900 ;
        RECT 25.240 13.840 25.450 14.165 ;
        RECT 8.990 13.680 11.530 13.840 ;
        RECT 8.390 13.560 11.530 13.680 ;
        RECT 23.960 13.630 25.450 13.840 ;
        RECT 8.390 13.400 9.270 13.560 ;
        RECT 23.960 13.480 24.190 13.630 ;
        RECT 1.680 13.140 2.000 13.170 ;
        RECT 2.660 13.140 2.890 13.335 ;
        RECT 1.680 12.940 2.890 13.140 ;
        RECT 1.680 12.910 2.000 12.940 ;
        RECT 2.660 12.795 2.890 12.940 ;
        RECT 8.990 12.360 9.270 13.400 ;
        RECT 23.695 13.290 23.985 13.320 ;
        RECT 24.380 13.290 25.345 13.345 ;
        RECT 23.695 13.115 25.345 13.290 ;
        RECT 23.695 13.090 23.985 13.115 ;
        RECT 25.115 13.005 25.345 13.115 ;
        RECT 26.715 13.005 26.945 14.165 ;
        RECT 29.690 13.290 34.460 13.520 ;
        RECT 29.690 13.005 29.920 13.290 ;
        RECT 34.095 13.280 34.385 13.290 ;
        RECT 25.115 12.775 29.920 13.005 ;
        RECT 10.180 12.670 10.460 12.700 ;
        RECT 10.180 12.390 11.600 12.670 ;
        RECT 29.690 12.495 29.920 12.775 ;
        RECT 34.095 12.495 34.385 12.540 ;
        RECT 10.180 12.360 10.460 12.390 ;
        RECT 29.690 12.265 34.455 12.495 ;
      LAYER met2 ;
        RECT 22.455 30.195 22.785 30.225 ;
        RECT 22.455 29.865 26.895 30.195 ;
        RECT 22.455 29.835 22.785 29.865 ;
        RECT 0.670 27.810 0.930 28.130 ;
        RECT 21.690 28.080 21.950 28.400 ;
        RECT 0.700 27.050 0.900 27.810 ;
        RECT 0.670 26.730 0.930 27.050 ;
        RECT 21.715 26.825 21.925 28.080 ;
        RECT 21.690 26.505 21.950 26.825 ;
        RECT 8.270 26.190 9.780 26.450 ;
        RECT -0.755 15.535 -0.345 15.885 ;
        RECT -3.750 15.365 -3.400 15.395 ;
        RECT -0.725 15.365 -0.375 15.535 ;
        RECT -3.750 15.015 -0.375 15.365 ;
        RECT -3.750 14.985 -3.400 15.015 ;
        RECT 1.710 13.980 1.970 14.300 ;
        RECT 1.740 13.200 1.940 13.980 ;
        RECT 1.710 12.880 1.970 13.200 ;
        RECT 8.960 12.390 10.490 12.670 ;
    END
  END VDD
  PIN down
    ANTENNAGATEAREA 2.872800 ;
    PORT
      LAYER li1 ;
        RECT 2.845 13.570 3.175 13.740 ;
        RECT 2.845 12.390 3.175 12.560 ;
        RECT 2.735 10.090 3.065 10.260 ;
        RECT 2.735 9.120 3.065 9.290 ;
        RECT 14.590 -0.105 14.760 0.225 ;
        RECT 30.140 -0.105 30.310 0.225 ;
      LAYER met1 ;
        RECT 2.865 13.760 3.155 13.770 ;
        RECT 0.640 13.550 3.170 13.760 ;
        RECT 0.640 12.515 0.850 13.550 ;
        RECT 2.865 13.540 3.155 13.550 ;
        RECT 2.865 12.515 3.155 12.590 ;
        RECT 0.640 12.305 3.195 12.515 ;
        RECT -1.240 11.600 -0.240 11.800 ;
        RECT 0.640 11.600 0.850 12.305 ;
        RECT -1.240 11.320 0.850 11.600 ;
        RECT -1.240 10.800 -0.240 11.320 ;
        RECT 0.030 4.740 0.310 11.320 ;
        RECT 0.640 10.255 0.850 11.320 ;
        RECT 2.755 10.255 3.045 10.290 ;
        RECT 0.640 10.045 3.095 10.255 ;
        RECT 0.640 9.265 0.850 10.045 ;
        RECT 2.755 9.265 3.045 9.320 ;
        RECT 0.640 9.090 3.045 9.265 ;
        RECT 0.640 9.055 3.025 9.090 ;
        RECT 3.700 4.740 3.975 4.770 ;
        RECT 7.980 4.740 8.255 4.770 ;
        RECT 0.030 4.460 2.630 4.740 ;
        RECT 3.700 4.465 7.195 4.740 ;
        RECT 7.980 4.465 18.835 4.740 ;
        RECT 3.700 4.435 3.975 4.465 ;
        RECT 7.980 4.435 8.255 4.465 ;
        RECT 14.580 1.665 14.770 1.700 ;
        RECT 18.560 1.665 18.835 4.465 ;
        RECT 14.580 1.475 30.265 1.665 ;
        RECT 14.580 0.205 14.770 1.475 ;
        RECT 18.560 1.415 18.835 1.475 ;
        RECT 30.075 0.205 30.265 1.475 ;
        RECT 14.560 -0.085 14.790 0.205 ;
        RECT 30.075 -0.035 30.340 0.205 ;
        RECT 30.110 -0.085 30.340 -0.035 ;
        RECT 14.580 -0.130 14.770 -0.085 ;
      LAYER met2 ;
        RECT 2.320 4.740 2.600 4.770 ;
        RECT 6.890 4.740 7.165 4.770 ;
        RECT 2.320 4.465 4.005 4.740 ;
        RECT 6.890 4.465 8.285 4.740 ;
        RECT 2.320 4.430 2.600 4.465 ;
        RECT 6.890 4.435 7.165 4.465 ;
    END
  END down
  PIN GND
    ANTENNAGATEAREA 0.345600 ;
    ANTENNADIFFAREA 14.725200 ;
    PORT
      LAYER pwell ;
        RECT 1.300 22.770 3.440 25.290 ;
        RECT 22.770 12.430 24.910 14.950 ;
        RECT 1.830 8.430 3.970 10.950 ;
        RECT 13.900 -1.010 31.000 1.130 ;
      LAYER li1 ;
        RECT 20.625 27.170 20.955 27.340 ;
        RECT 26.335 27.290 26.665 27.460 ;
        RECT 20.470 26.375 20.640 26.955 ;
        RECT 20.625 25.990 20.955 26.160 ;
        RECT 26.335 26.110 26.665 26.280 ;
        RECT 1.480 24.940 3.260 25.110 ;
        RECT 1.480 23.120 1.650 24.940 ;
        RECT 2.520 23.800 2.690 24.260 ;
        RECT 3.090 23.120 3.260 24.940 ;
        RECT 1.480 22.950 3.260 23.120 ;
        RECT 10.335 21.770 10.665 21.940 ;
        RECT 10.335 20.800 10.665 20.970 ;
        RECT 22.950 14.600 24.730 14.770 ;
        RECT 22.950 12.780 23.120 14.600 ;
        RECT 23.520 13.460 23.690 13.920 ;
        RECT 24.560 12.780 24.730 14.600 ;
        RECT 22.950 12.610 24.730 12.780 ;
        RECT 2.010 10.600 3.790 10.770 ;
        RECT 2.010 8.780 2.180 10.600 ;
        RECT 3.050 9.460 3.220 9.920 ;
        RECT 3.620 8.780 3.790 10.600 ;
        RECT 2.010 8.610 3.790 8.780 ;
        RECT 11.315 7.170 11.645 7.340 ;
        RECT 11.315 6.200 11.645 6.370 ;
        RECT 14.080 0.780 30.820 0.950 ;
        RECT 14.080 -0.660 14.250 0.780 ;
        RECT 14.930 -0.260 29.970 -0.090 ;
        RECT 30.650 -0.660 30.820 0.780 ;
        RECT 14.080 -0.830 30.820 -0.660 ;
      LAYER met1 ;
        RECT 68.640 87.180 73.450 87.700 ;
        RECT 68.640 72.900 69.160 87.180 ;
        RECT 68.610 71.900 73.350 72.900 ;
        RECT 68.640 66.760 69.160 71.900 ;
        RECT 77.810 71.870 78.810 72.930 ;
        RECT 68.610 66.240 69.190 66.760 ;
        RECT 68.640 47.480 69.160 62.450 ;
        RECT 64.260 46.960 69.160 47.480 ;
        RECT 20.640 27.150 22.540 27.400 ;
        RECT 20.645 27.140 20.935 27.150 ;
        RECT 20.440 26.720 20.670 26.935 ;
        RECT 19.340 26.520 20.670 26.720 ;
        RECT 2.490 24.210 2.720 24.240 ;
        RECT 2.490 23.960 3.770 24.210 ;
        RECT 19.340 23.970 19.540 26.520 ;
        RECT 20.440 26.395 20.670 26.520 ;
        RECT 22.290 26.825 22.540 27.150 ;
        RECT 24.550 27.270 26.670 27.510 ;
        RECT 24.550 26.825 24.790 27.270 ;
        RECT 26.355 27.260 26.645 27.270 ;
        RECT 22.290 26.575 24.790 26.825 ;
        RECT 22.290 26.280 22.540 26.575 ;
        RECT 24.550 26.320 24.790 26.575 ;
        RECT 24.550 26.310 26.640 26.320 ;
        RECT 22.290 26.245 22.570 26.280 ;
        RECT 20.655 26.190 22.570 26.245 ;
        RECT 20.645 25.995 22.570 26.190 ;
        RECT 24.550 26.080 26.645 26.310 ;
        RECT 20.645 25.960 20.935 25.995 ;
        RECT 22.370 23.970 22.570 25.995 ;
        RECT 2.490 23.820 2.720 23.960 ;
        RECT 3.520 23.195 3.770 23.960 ;
        RECT 2.605 23.150 3.770 23.195 ;
        RECT 1.510 22.945 3.770 23.150 ;
        RECT 14.920 23.770 22.570 23.970 ;
        RECT 1.510 22.480 3.370 22.945 ;
        RECT 2.240 16.750 2.520 22.480 ;
        RECT 7.700 22.000 7.980 22.030 ;
        RECT 6.850 21.720 7.980 22.000 ;
        RECT 8.790 21.720 10.680 22.000 ;
        RECT 6.850 21.020 7.130 21.720 ;
        RECT 7.700 21.690 7.980 21.720 ;
        RECT 6.850 20.740 10.690 21.020 ;
        RECT 6.850 16.750 7.130 20.740 ;
        RECT 14.920 19.070 15.120 23.770 ;
        RECT 14.890 18.750 15.150 19.070 ;
        RECT 14.860 17.080 15.180 17.340 ;
        RECT 14.920 16.750 15.120 17.080 ;
        RECT 2.210 16.705 15.280 16.750 ;
        RECT -1.945 16.395 15.280 16.705 ;
        RECT -1.945 3.470 -1.635 16.395 ;
        RECT 2.210 16.230 15.280 16.395 ;
        RECT 23.490 13.800 23.720 13.900 ;
        RECT 22.480 13.620 23.720 13.800 ;
        RECT 22.480 12.770 22.660 13.620 ;
        RECT 23.490 13.480 23.720 13.620 ;
        RECT 23.060 12.770 24.620 12.810 ;
        RECT 17.130 12.590 24.620 12.770 ;
        RECT 17.130 12.310 17.310 12.590 ;
        RECT 23.060 12.580 24.620 12.590 ;
        RECT 17.090 11.990 17.350 12.310 ;
        RECT 17.060 10.960 17.380 11.220 ;
        RECT 3.020 9.810 3.250 9.900 ;
        RECT 3.010 9.600 4.250 9.810 ;
        RECT 3.020 9.480 3.250 9.600 ;
        RECT 4.040 8.835 4.250 9.600 ;
        RECT 3.235 8.820 4.250 8.835 ;
        RECT 2.040 8.625 4.250 8.820 ;
        RECT 2.040 8.100 3.790 8.625 ;
        RECT 2.890 3.470 3.200 8.100 ;
        RECT 9.050 7.400 9.310 7.435 ;
        RECT 8.195 7.150 9.310 7.400 ;
        RECT 8.195 6.850 8.445 7.150 ;
        RECT 9.050 7.115 9.310 7.150 ;
        RECT 10.100 7.400 10.420 7.405 ;
        RECT 10.100 7.150 11.640 7.400 ;
        RECT 10.100 7.145 10.420 7.150 ;
        RECT 11.335 7.140 11.625 7.150 ;
        RECT 7.430 6.600 8.450 6.850 ;
        RECT 7.430 3.470 7.680 6.600 ;
        RECT 8.195 6.345 8.445 6.600 ;
        RECT 11.335 6.345 11.625 6.400 ;
        RECT 8.195 6.095 11.655 6.345 ;
        RECT 17.130 5.380 17.310 10.960 ;
        RECT 17.060 5.120 17.380 5.380 ;
        RECT 17.060 3.840 17.380 4.100 ;
        RECT -1.945 3.420 16.930 3.470 ;
        RECT 17.130 3.420 17.310 3.840 ;
        RECT -1.945 3.170 17.440 3.420 ;
        RECT -1.945 3.160 8.970 3.170 ;
        RECT 11.090 3.160 17.440 3.170 ;
        RECT 6.830 -4.750 7.270 3.160 ;
        RECT 13.605 0.840 13.915 3.160 ;
        RECT 13.605 0.495 14.280 0.840 ;
        RECT 13.700 -0.800 14.280 0.495 ;
        RECT 15.280 -0.060 15.480 -0.030 ;
        RECT 15.035 -0.290 21.105 -0.060 ;
        RECT 14.010 -1.160 14.210 -0.800 ;
        RECT 15.280 -1.160 15.480 -0.290 ;
        RECT 14.010 -1.360 15.480 -1.160 ;
        RECT 78.090 -4.750 78.530 71.870 ;
        RECT 6.830 -5.190 78.530 -4.750 ;
      LAYER met2 ;
        RECT 72.900 87.700 73.420 87.730 ;
        RECT 72.900 87.180 77.705 87.700 ;
        RECT 72.900 87.150 73.420 87.180 ;
        RECT 72.320 72.900 73.320 72.930 ;
        RECT 72.320 71.900 78.840 72.900 ;
        RECT 72.320 71.870 73.320 71.900 ;
        RECT 68.640 62.420 69.160 66.790 ;
        RECT 68.610 61.900 69.190 62.420 ;
        RECT 64.290 47.480 64.810 47.510 ;
        RECT 62.365 46.960 64.810 47.480 ;
        RECT 64.290 46.930 64.810 46.960 ;
        RECT 8.820 22.000 9.100 22.030 ;
        RECT 7.670 21.720 9.100 22.000 ;
        RECT 8.820 21.690 9.100 21.720 ;
        RECT 14.860 18.780 15.180 19.040 ;
        RECT 14.920 17.370 15.120 18.780 ;
        RECT 14.890 17.050 15.150 17.370 ;
        RECT 17.060 12.020 17.380 12.280 ;
        RECT 17.130 11.250 17.310 12.020 ;
        RECT 17.090 10.930 17.350 11.250 ;
        RECT 9.020 7.400 9.340 7.405 ;
        RECT 10.130 7.400 10.390 7.435 ;
        RECT 9.020 7.150 10.390 7.400 ;
        RECT 9.020 7.145 9.340 7.150 ;
        RECT 10.130 7.115 10.390 7.150 ;
        RECT 17.090 5.090 17.350 5.410 ;
        RECT 17.130 4.130 17.310 5.090 ;
        RECT 17.090 3.810 17.350 4.130 ;
      LAYER met3 ;
        RECT -322.220 410.650 -291.820 442.510 ;
        RECT -290.620 410.650 -260.220 442.510 ;
        RECT -259.020 410.650 -228.620 442.510 ;
        RECT -227.420 410.650 -197.020 442.510 ;
        RECT -195.820 410.650 -165.420 442.510 ;
        RECT -164.220 410.650 -133.820 442.510 ;
        RECT -132.620 410.650 -102.220 442.510 ;
        RECT -101.020 410.650 -70.620 442.510 ;
        RECT -69.420 410.650 -39.020 442.510 ;
        RECT -37.820 410.650 -7.420 442.510 ;
        RECT -6.220 410.650 24.180 442.510 ;
        RECT 25.380 410.650 55.780 442.510 ;
        RECT -324.780 392.785 -324.260 395.750 ;
        RECT -324.805 392.275 -324.235 392.785 ;
        RECT -324.780 392.270 -324.260 392.275 ;
        RECT -322.220 377.590 -291.820 409.450 ;
        RECT -290.620 377.590 -260.220 409.450 ;
        RECT -259.020 377.590 -228.620 409.450 ;
        RECT -227.420 377.590 -197.020 409.450 ;
        RECT -195.820 377.590 -165.420 409.450 ;
        RECT -164.220 377.590 -133.820 409.450 ;
        RECT -132.620 377.590 -102.220 409.450 ;
        RECT -101.020 377.590 -70.620 409.450 ;
        RECT -69.420 377.590 -39.020 409.450 ;
        RECT -37.820 377.590 -7.420 409.450 ;
        RECT -6.220 377.590 24.180 409.450 ;
        RECT 25.380 377.590 55.780 409.450 ;
        RECT -322.220 344.530 -291.820 376.390 ;
        RECT -290.620 344.530 -260.220 376.390 ;
        RECT -259.020 344.530 -228.620 376.390 ;
        RECT -227.420 344.530 -197.020 376.390 ;
        RECT -195.820 344.530 -165.420 376.390 ;
        RECT -164.220 344.530 -133.820 376.390 ;
        RECT -132.620 344.530 -102.220 376.390 ;
        RECT -101.020 344.530 -70.620 376.390 ;
        RECT -69.420 344.530 -39.020 376.390 ;
        RECT -37.820 344.530 -7.420 376.390 ;
        RECT -6.220 344.530 24.180 376.390 ;
        RECT 25.380 344.530 55.780 376.390 ;
        RECT 56.800 359.210 57.320 362.780 ;
        RECT 56.805 359.185 57.315 359.210 ;
        RECT -323.910 327.005 -323.390 329.280 ;
        RECT -323.935 326.495 -323.365 327.005 ;
        RECT -323.910 326.490 -323.390 326.495 ;
        RECT -322.220 311.470 -291.820 343.330 ;
        RECT -290.620 311.470 -260.220 343.330 ;
        RECT -259.020 311.470 -228.620 343.330 ;
        RECT -227.420 311.470 -197.020 343.330 ;
        RECT -195.820 311.470 -165.420 343.330 ;
        RECT -164.220 311.470 -133.820 343.330 ;
        RECT -132.620 311.470 -102.220 343.330 ;
        RECT -101.020 311.470 -70.620 343.330 ;
        RECT -69.420 311.470 -39.020 343.330 ;
        RECT -37.820 311.470 -7.420 343.330 ;
        RECT -6.220 311.470 24.180 343.330 ;
        RECT 25.380 311.470 55.780 343.330 ;
        RECT -322.220 278.410 -291.820 310.270 ;
        RECT -290.620 278.410 -260.220 310.270 ;
        RECT -259.020 278.410 -228.620 310.270 ;
        RECT -227.420 278.410 -197.020 310.270 ;
        RECT -195.820 278.410 -165.420 310.270 ;
        RECT -164.220 278.410 -133.820 310.270 ;
        RECT -132.620 278.410 -102.220 310.270 ;
        RECT -101.020 278.410 -70.620 310.270 ;
        RECT -69.420 278.410 -39.020 310.270 ;
        RECT -37.820 278.410 -7.420 310.270 ;
        RECT -6.220 278.410 24.180 310.270 ;
        RECT 25.380 278.410 55.780 310.270 ;
        RECT 56.850 293.925 57.370 297.260 ;
        RECT 56.825 293.415 57.395 293.925 ;
        RECT 56.850 293.410 57.370 293.415 ;
        RECT -324.060 260.875 -323.540 263.300 ;
        RECT -324.085 260.365 -323.515 260.875 ;
        RECT -324.060 260.360 -323.540 260.365 ;
        RECT -322.220 245.350 -291.820 277.210 ;
        RECT -290.620 245.350 -260.220 277.210 ;
        RECT -259.020 245.350 -228.620 277.210 ;
        RECT -227.420 245.350 -197.020 277.210 ;
        RECT -195.820 245.350 -165.420 277.210 ;
        RECT -164.220 245.350 -133.820 277.210 ;
        RECT -132.620 245.350 -102.220 277.210 ;
        RECT -101.020 245.350 -70.620 277.210 ;
        RECT -69.420 245.350 -39.020 277.210 ;
        RECT -37.820 245.350 -7.420 277.210 ;
        RECT -6.220 245.350 24.180 277.210 ;
        RECT 25.380 245.350 55.780 277.210 ;
        RECT -322.220 212.290 -291.820 244.150 ;
        RECT -290.620 212.290 -260.220 244.150 ;
        RECT -259.020 212.290 -228.620 244.150 ;
        RECT -227.420 212.290 -197.020 244.150 ;
        RECT -195.820 212.290 -165.420 244.150 ;
        RECT -164.220 212.290 -133.820 244.150 ;
        RECT -132.620 212.290 -102.220 244.150 ;
        RECT -101.020 212.290 -70.620 244.150 ;
        RECT -69.420 212.290 -39.020 244.150 ;
        RECT -37.820 212.290 -7.420 244.150 ;
        RECT -6.220 212.290 24.180 244.150 ;
        RECT 25.380 212.290 55.780 244.150 ;
        RECT 56.890 227.685 57.410 230.450 ;
        RECT 56.865 227.175 57.435 227.685 ;
        RECT 56.890 227.170 57.410 227.175 ;
        RECT 92.755 214.320 96.625 214.325 ;
        RECT 92.730 213.795 96.625 214.320 ;
        RECT 97.830 213.800 128.230 245.660 ;
        RECT 129.430 213.800 159.830 245.660 ;
        RECT 161.030 213.800 191.430 245.660 ;
        RECT 192.630 213.800 223.030 245.660 ;
        RECT 224.230 213.800 254.630 245.660 ;
        RECT 92.755 213.790 96.625 213.795 ;
        RECT -324.460 194.290 -323.940 197.380 ;
        RECT -324.455 194.265 -323.945 194.290 ;
        RECT -322.220 179.230 -291.820 211.090 ;
        RECT -290.620 179.230 -260.220 211.090 ;
        RECT -259.020 179.230 -228.620 211.090 ;
        RECT -227.420 179.230 -197.020 211.090 ;
        RECT -195.820 179.230 -165.420 211.090 ;
        RECT -164.220 179.230 -133.820 211.090 ;
        RECT -132.620 179.230 -102.220 211.090 ;
        RECT -101.020 179.230 -70.620 211.090 ;
        RECT -69.420 179.230 -39.020 211.090 ;
        RECT -37.820 179.230 -7.420 211.090 ;
        RECT -6.220 179.230 24.180 211.090 ;
        RECT 25.380 179.230 55.780 211.090 ;
        RECT 97.830 180.740 128.230 212.600 ;
        RECT 129.430 180.740 159.830 212.600 ;
        RECT 161.030 180.740 191.430 212.600 ;
        RECT 192.630 180.740 223.030 212.600 ;
        RECT 224.230 180.740 254.630 212.600 ;
        RECT -322.220 146.170 -291.820 178.030 ;
        RECT -290.620 146.170 -260.220 178.030 ;
        RECT -259.020 146.170 -228.620 178.030 ;
        RECT -227.420 146.170 -197.020 178.030 ;
        RECT -195.820 146.170 -165.420 178.030 ;
        RECT -164.220 146.170 -133.820 178.030 ;
        RECT -132.620 146.170 -102.220 178.030 ;
        RECT -101.020 146.170 -70.620 178.030 ;
        RECT -69.420 146.170 -39.020 178.030 ;
        RECT -37.820 146.170 -7.420 178.030 ;
        RECT -6.220 146.170 24.180 178.030 ;
        RECT 25.380 146.170 55.780 178.030 ;
        RECT 57.080 161.765 57.600 164.340 ;
        RECT 57.055 161.255 57.625 161.765 ;
        RECT 57.080 161.250 57.600 161.255 ;
        RECT 97.830 147.680 128.230 179.540 ;
        RECT 129.430 147.680 159.830 179.540 ;
        RECT 161.030 147.680 191.430 179.540 ;
        RECT 192.630 147.680 223.030 179.540 ;
        RECT 224.230 147.680 254.630 179.540 ;
        RECT -324.240 128.735 -323.720 131.250 ;
        RECT -324.265 128.225 -323.695 128.735 ;
        RECT -324.240 128.220 -323.720 128.225 ;
        RECT -322.220 113.110 -291.820 144.970 ;
        RECT -290.620 113.110 -260.220 144.970 ;
        RECT -259.020 113.110 -228.620 144.970 ;
        RECT -227.420 113.110 -197.020 144.970 ;
        RECT -195.820 113.110 -165.420 144.970 ;
        RECT -164.220 113.110 -133.820 144.970 ;
        RECT -132.620 113.110 -102.220 144.970 ;
        RECT -101.020 113.110 -70.620 144.970 ;
        RECT -69.420 113.110 -39.020 144.970 ;
        RECT -37.820 113.110 -7.420 144.970 ;
        RECT -6.220 113.110 24.180 144.970 ;
        RECT 25.380 113.110 55.780 144.970 ;
        RECT 95.640 129.975 96.160 133.080 ;
        RECT 95.615 129.465 96.185 129.975 ;
        RECT 95.640 129.460 96.160 129.465 ;
        RECT 97.830 114.620 128.230 146.480 ;
        RECT 129.430 114.620 159.830 146.480 ;
        RECT 161.030 114.620 191.430 146.480 ;
        RECT 192.630 114.620 223.030 146.480 ;
        RECT 224.230 114.620 254.630 146.480 ;
        RECT 255.600 115.155 258.810 115.160 ;
        RECT 255.600 114.645 258.835 115.155 ;
        RECT 255.600 114.640 258.810 114.645 ;
        RECT -322.220 80.050 -291.820 111.910 ;
        RECT -290.620 80.050 -260.220 111.910 ;
        RECT -259.020 80.050 -228.620 111.910 ;
        RECT -227.420 80.050 -197.020 111.910 ;
        RECT -195.820 80.050 -165.420 111.910 ;
        RECT -164.220 80.050 -133.820 111.910 ;
        RECT -132.620 80.050 -102.220 111.910 ;
        RECT -101.020 80.050 -70.620 111.910 ;
        RECT -69.420 80.050 -39.020 111.910 ;
        RECT -37.820 80.050 -7.420 111.910 ;
        RECT -6.220 80.050 24.180 111.910 ;
        RECT 25.380 80.050 55.780 111.910 ;
        RECT 57.120 95.695 57.640 98.050 ;
        RECT 57.095 95.185 57.665 95.695 ;
        RECT 57.120 95.180 57.640 95.185 ;
        RECT 77.115 87.700 77.685 87.725 ;
        RECT 77.115 87.180 83.470 87.700 ;
        RECT 77.115 87.155 77.685 87.180 ;
        RECT 97.830 81.560 128.230 113.420 ;
        RECT 129.430 81.560 159.830 113.420 ;
        RECT 161.030 81.560 191.430 113.420 ;
        RECT 192.630 81.560 223.030 113.420 ;
        RECT 224.230 81.560 254.630 113.420 ;
        RECT -325.110 62.395 -324.590 66.000 ;
        RECT -325.135 61.885 -324.565 62.395 ;
        RECT -325.110 61.880 -324.590 61.885 ;
        RECT -322.220 46.990 -291.820 78.850 ;
        RECT -290.620 46.990 -260.220 78.850 ;
        RECT -259.020 46.990 -228.620 78.850 ;
        RECT -227.420 46.990 -197.020 78.850 ;
        RECT -195.820 46.990 -165.420 78.850 ;
        RECT -164.220 46.990 -133.820 78.850 ;
        RECT -132.620 46.990 -102.220 78.850 ;
        RECT -101.020 46.990 -70.620 78.850 ;
        RECT -69.420 46.990 -39.020 78.850 ;
        RECT -37.820 46.990 -7.420 78.850 ;
        RECT -6.220 46.990 24.180 78.850 ;
        RECT 25.380 46.990 55.780 78.850 ;
        RECT 62.385 47.480 62.955 47.505 ;
        RECT 59.890 46.960 62.955 47.480 ;
        RECT 62.385 46.935 62.955 46.960 ;
      LAYER met4 ;
        RECT -322.820 411.110 56.380 411.170 ;
        RECT -324.780 410.650 56.380 411.110 ;
        RECT -324.780 410.590 -322.380 410.650 ;
        RECT -324.780 395.725 -324.260 410.590 ;
        RECT -324.785 395.195 -324.255 395.725 ;
        RECT -324.780 378.110 -324.260 392.790 ;
        RECT -324.780 378.085 56.380 378.110 ;
        RECT -324.780 377.590 57.325 378.085 ;
        RECT 55.915 377.555 57.325 377.590 ;
        RECT 56.795 362.225 57.325 377.555 ;
        RECT 56.800 345.050 57.320 359.730 ;
        RECT -322.820 345.010 57.320 345.050 ;
        RECT -323.910 344.530 57.320 345.010 ;
        RECT -323.910 344.490 -322.230 344.530 ;
        RECT -323.910 329.255 -323.390 344.490 ;
        RECT -323.915 328.725 -323.385 329.255 ;
        RECT -323.910 311.990 -323.390 327.010 ;
        RECT 55.810 311.990 57.370 312.040 ;
        RECT -323.910 311.520 57.370 311.990 ;
        RECT -323.910 311.470 56.380 311.520 ;
        RECT 56.850 297.235 57.370 311.520 ;
        RECT 56.845 296.705 57.375 297.235 ;
        RECT 56.850 278.930 57.370 293.930 ;
        RECT -322.820 278.830 57.370 278.930 ;
        RECT -324.060 278.410 57.370 278.830 ;
        RECT -324.060 278.310 -322.410 278.410 ;
        RECT -324.060 263.275 -323.540 278.310 ;
        RECT -324.065 262.745 -323.535 263.275 ;
        RECT -324.060 245.870 -323.540 260.880 ;
        RECT 56.040 245.870 57.410 245.910 ;
        RECT -324.060 245.390 57.410 245.870 ;
        RECT -324.060 245.350 56.380 245.390 ;
        RECT 56.890 230.425 57.410 245.390 ;
        RECT 56.885 229.895 57.415 230.425 ;
        RECT -324.460 212.810 -321.900 212.840 ;
        RECT 56.890 212.810 57.410 227.690 ;
        RECT 96.055 214.325 96.600 214.330 ;
        RECT -324.460 212.320 57.410 212.810 ;
        RECT -324.460 197.355 -323.940 212.320 ;
        RECT -322.820 212.290 57.410 212.320 ;
        RECT -324.465 196.825 -323.935 197.355 ;
        RECT -324.460 179.750 -323.940 194.810 ;
        RECT 92.755 181.260 93.290 214.325 ;
        RECT 96.055 214.320 97.695 214.325 ;
        RECT 96.055 213.800 255.230 214.320 ;
        RECT 96.055 213.790 97.695 213.800 ;
        RECT 96.055 213.785 96.600 213.790 ;
        RECT 254.935 181.260 258.440 181.265 ;
        RECT 92.755 180.750 258.440 181.260 ;
        RECT 92.755 180.740 255.230 180.750 ;
        RECT 92.755 180.735 93.290 180.740 ;
        RECT -324.460 179.690 56.380 179.750 ;
        RECT -324.460 179.230 57.600 179.690 ;
        RECT 56.170 179.170 57.600 179.230 ;
        RECT 57.080 164.315 57.600 179.170 ;
        RECT 57.075 163.785 57.605 164.315 ;
        RECT -324.240 146.690 -322.400 146.720 ;
        RECT 57.080 146.690 57.600 161.770 ;
        RECT 257.925 148.200 258.440 180.750 ;
        RECT 97.230 148.150 258.440 148.200 ;
        RECT -324.240 146.200 57.600 146.690 ;
        RECT -324.240 131.225 -323.720 146.200 ;
        RECT -322.820 146.170 57.600 146.200 ;
        RECT 95.640 147.680 258.440 148.150 ;
        RECT 95.640 147.630 97.560 147.680 ;
        RECT 95.640 133.055 96.160 147.630 ;
        RECT 95.635 132.525 96.165 133.055 ;
        RECT -324.245 130.695 -323.715 131.225 ;
        RECT -324.240 113.630 -323.720 128.740 ;
        RECT 95.640 115.140 96.160 129.980 ;
        RECT 255.625 115.160 256.155 115.165 ;
        RECT 254.680 115.140 256.155 115.160 ;
        RECT 95.640 114.640 256.155 115.140 ;
        RECT 95.640 114.620 255.230 114.640 ;
        RECT 255.625 114.635 256.155 114.640 ;
        RECT 55.930 113.630 57.640 113.720 ;
        RECT -324.240 113.200 57.640 113.630 ;
        RECT -324.240 113.110 56.380 113.200 ;
        RECT 57.120 98.025 57.640 113.200 ;
        RECT 57.115 97.495 57.645 98.025 ;
        RECT -325.110 80.570 -322.190 80.620 ;
        RECT 57.120 80.570 57.640 95.700 ;
        RECT 82.915 87.700 83.445 87.705 ;
        RECT 82.915 87.180 96.130 87.700 ;
        RECT 82.915 87.175 83.445 87.180 ;
        RECT 95.610 82.060 96.130 87.180 ;
        RECT 258.290 82.080 258.810 115.160 ;
        RECT 97.230 82.060 258.810 82.080 ;
        RECT 95.610 81.560 258.810 82.060 ;
        RECT 95.610 81.540 97.680 81.560 ;
        RECT -325.110 80.100 57.640 80.570 ;
        RECT -325.110 65.975 -324.590 80.100 ;
        RECT -322.820 80.050 57.640 80.100 ;
        RECT -325.115 65.445 -324.585 65.975 ;
        RECT -325.110 47.510 -324.590 62.400 ;
        RECT -325.110 47.480 57.400 47.510 ;
        RECT 59.915 47.480 60.445 47.485 ;
        RECT -325.110 46.990 60.445 47.480 ;
        RECT 56.830 46.960 60.445 46.990 ;
        RECT 59.915 46.955 60.445 46.960 ;
    END
  END GND
  OBS
      LAYER pwell ;
        RECT 56.690 36.070 58.830 43.680 ;
      LAYER nwell ;
        RECT 9.410 24.090 11.550 28.280 ;
        RECT 25.430 25.420 27.570 28.150 ;
        RECT 9.350 24.080 11.550 24.090 ;
        RECT 7.600 22.650 13.410 24.080 ;
        RECT 7.600 20.080 9.030 22.650 ;
      LAYER pwell ;
        RECT 9.430 20.110 11.570 22.630 ;
      LAYER nwell ;
        RECT 11.980 20.080 13.410 22.650 ;
        RECT 7.600 18.650 13.410 20.080 ;
        RECT 17.540 17.930 19.680 20.660 ;
        RECT 10.300 9.500 12.440 14.500 ;
        RECT 31.310 14.180 37.120 15.610 ;
        RECT 31.310 11.610 32.740 14.180 ;
      LAYER pwell ;
        RECT 33.170 11.650 35.310 14.170 ;
      LAYER nwell ;
        RECT 35.690 11.610 37.120 14.180 ;
        RECT 8.660 8.070 14.470 9.500 ;
        RECT 8.660 5.500 10.090 8.070 ;
      LAYER pwell ;
        RECT 10.410 5.510 12.550 8.030 ;
      LAYER nwell ;
        RECT 13.040 5.500 14.470 8.070 ;
        RECT 8.660 4.070 14.470 5.500 ;
        RECT 19.980 9.380 25.790 10.810 ;
        RECT 31.310 10.180 37.120 11.610 ;
        RECT 19.980 6.810 21.410 9.380 ;
      LAYER pwell ;
        RECT 21.870 6.820 24.010 9.340 ;
      LAYER nwell ;
        RECT 24.360 6.810 25.790 9.380 ;
        RECT 19.980 5.380 25.790 6.810 ;
      LAYER li1 ;
        RECT 56.870 43.330 58.650 43.500 ;
        RECT 56.870 36.420 57.040 43.330 ;
        RECT 57.520 42.600 58.000 42.770 ;
        RECT 57.600 40.785 57.920 42.600 ;
        RECT 58.480 36.420 58.650 43.330 ;
        RECT 56.870 36.250 58.650 36.420 ;
        RECT -5.100 32.935 -4.930 33.265 ;
        RECT -4.715 32.780 40.325 32.950 ;
        RECT 40.540 32.935 40.710 33.265 ;
        RECT 9.590 27.930 11.370 28.100 ;
        RECT 2.500 26.575 2.670 27.155 ;
        RECT 9.590 25.900 9.760 27.930 ;
        RECT 10.160 26.625 10.330 27.205 ;
        RECT 10.630 26.625 10.800 27.205 ;
        RECT 11.200 25.900 11.370 27.930 ;
        RECT 9.590 25.730 11.370 25.900 ;
        RECT 25.610 27.800 27.390 27.970 ;
        RECT 25.610 25.770 25.780 27.800 ;
        RECT 26.180 26.495 26.350 27.075 ;
        RECT 27.220 25.770 27.390 27.800 ;
        RECT 25.610 25.600 27.390 25.770 ;
        RECT 2.050 23.800 2.220 24.260 ;
        RECT 7.885 23.625 13.125 23.795 ;
        RECT 7.885 19.105 8.055 23.625 ;
        RECT 9.610 22.280 11.390 22.450 ;
        RECT 9.610 20.460 9.780 22.280 ;
        RECT 10.180 21.140 10.350 21.600 ;
        RECT 10.650 21.140 10.820 21.600 ;
        RECT 11.220 20.460 11.390 22.280 ;
        RECT 9.610 20.290 11.390 20.460 ;
        RECT 12.955 19.105 13.125 23.625 ;
        RECT 7.885 18.935 13.125 19.105 ;
        RECT 17.720 20.310 19.500 20.480 ;
        RECT 17.720 18.280 17.890 20.310 ;
        RECT 18.290 19.005 18.460 19.585 ;
        RECT 18.760 19.005 18.930 19.585 ;
        RECT 19.330 18.280 19.500 20.310 ;
        RECT 17.720 18.110 19.500 18.280 ;
        RECT 31.595 15.155 36.835 15.325 ;
        RECT 10.480 14.150 12.260 14.320 ;
        RECT 3.160 12.775 3.330 13.355 ;
        RECT 10.480 12.120 10.650 14.150 ;
        RECT 11.050 12.845 11.220 13.425 ;
        RECT 11.520 12.845 11.690 13.425 ;
        RECT 12.090 12.120 12.260 14.150 ;
        RECT 10.480 11.950 12.260 12.120 ;
        RECT 31.595 10.635 31.765 15.155 ;
        RECT 33.350 13.820 35.130 13.990 ;
        RECT 33.350 12.000 33.520 13.820 ;
        RECT 34.390 12.680 34.560 13.140 ;
        RECT 34.960 12.000 35.130 13.820 ;
        RECT 33.350 11.830 35.130 12.000 ;
        RECT 36.665 10.635 36.835 15.155 ;
        RECT 20.265 10.355 25.505 10.525 ;
        RECT 31.595 10.465 36.835 10.635 ;
        RECT 2.580 9.460 2.750 9.920 ;
        RECT 8.945 9.045 14.185 9.215 ;
        RECT 8.945 4.525 9.115 9.045 ;
        RECT 10.590 7.680 12.370 7.850 ;
        RECT 10.590 5.860 10.760 7.680 ;
        RECT 11.160 6.540 11.330 7.000 ;
        RECT 11.630 6.540 11.800 7.000 ;
        RECT 12.200 5.860 12.370 7.680 ;
        RECT 10.590 5.690 12.370 5.860 ;
        RECT 14.015 4.525 14.185 9.045 ;
        RECT 20.265 5.835 20.435 10.355 ;
        RECT 22.050 8.990 23.830 9.160 ;
        RECT 22.050 7.170 22.220 8.990 ;
        RECT 22.775 8.480 23.105 8.650 ;
        RECT 22.620 7.850 22.790 8.310 ;
        RECT 23.090 7.850 23.260 8.310 ;
        RECT 22.775 7.510 23.105 7.680 ;
        RECT 23.660 7.170 23.830 8.990 ;
        RECT 22.050 7.000 23.830 7.170 ;
        RECT 25.335 5.835 25.505 10.355 ;
        RECT 20.265 5.665 25.505 5.835 ;
        RECT 8.945 4.355 14.185 4.525 ;
        RECT 14.930 0.210 29.970 0.380 ;
      LAYER met1 ;
        RECT 61.550 63.910 62.070 63.940 ;
        RECT 61.550 63.390 72.770 63.910 ;
        RECT 61.550 63.360 62.070 63.390 ;
        RECT 72.250 45.450 72.770 63.390 ;
        RECT 57.560 44.930 72.770 45.450 ;
        RECT 57.560 43.730 58.080 44.930 ;
        RECT 57.600 42.830 57.920 43.730 ;
        RECT 57.570 40.725 57.950 42.830 ;
        RECT -5.180 31.900 -4.900 33.280 ;
        RECT -4.610 32.750 13.460 32.980 ;
        RECT 12.110 32.100 12.370 32.750 ;
        RECT 13.870 31.900 14.030 31.920 ;
        RECT 40.480 31.900 40.760 33.250 ;
        RECT -5.180 31.620 40.760 31.900 ;
        RECT 12.080 31.050 13.670 31.310 ;
        RECT 13.870 29.590 14.030 31.620 ;
        RECT 14.660 31.310 14.920 31.340 ;
        RECT 14.660 31.050 25.920 31.310 ;
        RECT 14.660 31.020 14.920 31.050 ;
        RECT 13.790 29.330 14.110 29.590 ;
        RECT 13.820 27.720 14.080 28.040 ;
        RECT 23.695 27.970 23.925 31.050 ;
        RECT 25.740 28.550 25.920 31.050 ;
        RECT 25.740 28.370 26.610 28.550 ;
        RECT 25.740 28.180 25.920 28.370 ;
        RECT 2.470 26.960 2.700 27.135 ;
        RECT 10.130 27.000 10.360 27.185 ;
        RECT 2.470 26.740 3.740 26.960 ;
        RECT 2.470 26.595 2.700 26.740 ;
        RECT 1.100 25.500 1.420 25.520 ;
        RECT 3.520 25.500 3.740 26.740 ;
        RECT 9.090 26.840 10.360 27.000 ;
        RECT 9.090 25.590 9.250 26.840 ;
        RECT 10.130 26.645 10.360 26.840 ;
        RECT 10.600 27.060 10.830 27.185 ;
        RECT 10.600 26.850 11.990 27.060 ;
        RECT 10.600 26.645 10.830 26.850 ;
        RECT 9.700 25.830 11.260 25.930 ;
        RECT 9.500 25.640 11.390 25.830 ;
        RECT 9.500 25.590 11.540 25.640 ;
        RECT 1.100 25.280 6.840 25.500 ;
        RECT 9.090 25.430 11.540 25.590 ;
        RECT 11.220 25.380 11.540 25.430 ;
        RECT 1.100 25.260 1.420 25.280 ;
        RECT 6.620 24.480 6.840 25.280 ;
        RECT 11.780 24.525 11.990 26.850 ;
        RECT 12.440 25.350 12.700 25.670 ;
        RECT 8.355 24.480 11.990 24.525 ;
        RECT 6.620 24.315 11.990 24.480 ;
        RECT 12.490 24.680 12.650 25.350 ;
        RECT 13.870 24.680 14.030 27.720 ;
        RECT 23.680 27.650 23.940 27.970 ;
        RECT 25.700 27.860 25.960 28.180 ;
        RECT 26.430 28.010 26.610 28.370 ;
        RECT 26.300 28.000 27.220 28.010 ;
        RECT 26.300 27.800 27.280 28.000 ;
        RECT 26.585 27.770 27.280 27.800 ;
        RECT 25.670 26.850 25.990 26.890 ;
        RECT 26.150 26.850 26.380 27.055 ;
        RECT 25.670 26.670 26.380 26.850 ;
        RECT 25.670 26.630 25.990 26.670 ;
        RECT 26.150 26.515 26.380 26.670 ;
        RECT 23.680 25.740 23.940 26.060 ;
        RECT 12.490 24.520 14.030 24.680 ;
        RECT 6.620 24.260 8.565 24.315 ;
        RECT 1.100 24.110 1.420 24.130 ;
        RECT 2.020 24.110 2.250 24.240 ;
        RECT 1.100 23.890 2.250 24.110 ;
        RECT 1.100 23.870 1.420 23.890 ;
        RECT 2.020 23.820 2.250 23.890 ;
        RECT 8.355 21.445 8.565 24.260 ;
        RECT 10.150 21.445 10.380 21.580 ;
        RECT 8.355 21.235 10.380 21.445 ;
        RECT 10.150 21.160 10.380 21.235 ;
        RECT 10.620 21.390 10.850 21.580 ;
        RECT 12.490 21.390 12.650 24.520 ;
        RECT 10.620 21.230 12.650 21.390 ;
        RECT 10.620 21.160 10.850 21.230 ;
        RECT 9.720 20.470 11.280 20.490 ;
        RECT 11.790 20.470 11.950 21.230 ;
        RECT 9.720 20.310 11.950 20.470 ;
        RECT 9.720 20.260 11.280 20.310 ;
        RECT 18.260 19.460 18.490 19.565 ;
        RECT 18.730 19.460 18.960 19.565 ;
        RECT 19.300 19.460 19.530 20.370 ;
        RECT 23.695 19.460 23.925 25.740 ;
        RECT 18.260 19.230 23.925 19.460 ;
        RECT 18.260 19.025 18.490 19.230 ;
        RECT 18.730 19.025 18.960 19.230 ;
        RECT 19.300 18.220 19.530 19.230 ;
        RECT 3.130 13.140 3.360 13.335 ;
        RECT 11.020 13.150 11.250 13.405 ;
        RECT 3.130 12.950 4.470 13.140 ;
        RECT 3.130 12.795 3.360 12.950 ;
        RECT 4.280 11.760 4.470 12.950 ;
        RECT 9.840 12.970 11.250 13.150 ;
        RECT 9.840 11.810 10.020 12.970 ;
        RECT 11.020 12.865 11.250 12.970 ;
        RECT 11.490 13.250 11.720 13.405 ;
        RECT 11.490 13.080 13.050 13.250 ;
        RECT 11.490 12.865 11.720 13.080 ;
        RECT 10.590 12.000 12.150 12.150 ;
        RECT 10.420 11.980 12.260 12.000 ;
        RECT 10.420 11.850 12.360 11.980 ;
        RECT 10.420 11.810 12.620 11.850 ;
        RECT 4.280 11.480 8.400 11.760 ;
        RECT 9.840 11.630 12.620 11.810 ;
        RECT 4.280 11.325 4.470 11.480 ;
        RECT 1.935 11.135 4.470 11.325 ;
        RECT 1.935 10.930 2.125 11.135 ;
        RECT 1.900 10.610 2.160 10.930 ;
        RECT 8.120 10.245 8.400 11.480 ;
        RECT 12.270 11.590 12.620 11.630 ;
        RECT 12.270 10.680 12.450 11.590 ;
        RECT 12.230 10.360 12.490 10.680 ;
        RECT 8.120 10.195 10.030 10.245 ;
        RECT 12.880 10.195 13.050 13.080 ;
        RECT 34.360 13.065 34.590 13.120 ;
        RECT 34.360 12.875 35.535 13.065 ;
        RECT 34.360 12.700 34.590 12.875 ;
        RECT 33.460 11.985 35.020 12.030 ;
        RECT 35.345 11.985 35.535 12.875 ;
        RECT 13.280 11.810 13.540 11.880 ;
        RECT 13.280 11.630 19.230 11.810 ;
        RECT 33.460 11.800 35.535 11.985 ;
        RECT 13.280 11.560 13.540 11.630 ;
        RECT 8.120 10.080 13.050 10.195 ;
        RECT 8.120 10.020 8.400 10.080 ;
        RECT 9.585 10.025 13.050 10.080 ;
        RECT 1.870 9.805 2.190 9.840 ;
        RECT 2.550 9.805 2.780 9.900 ;
        RECT 1.870 9.615 2.780 9.805 ;
        RECT 1.870 9.580 2.190 9.615 ;
        RECT 2.550 9.480 2.780 9.615 ;
        RECT 9.585 6.775 9.755 10.025 ;
        RECT 12.200 9.420 12.520 9.680 ;
        RECT 11.130 6.775 11.360 6.980 ;
        RECT 9.585 6.605 11.360 6.775 ;
        RECT 11.130 6.560 11.360 6.605 ;
        RECT 11.600 6.810 11.830 6.980 ;
        RECT 12.270 6.810 12.450 9.420 ;
        RECT 19.050 8.110 19.230 11.630 ;
        RECT 34.715 11.795 35.535 11.800 ;
        RECT 22.070 8.510 23.100 8.690 ;
        RECT 22.070 8.110 22.250 8.510 ;
        RECT 22.795 8.450 23.085 8.510 ;
        RECT 22.590 8.190 22.820 8.290 ;
        RECT 23.060 8.190 23.290 8.290 ;
        RECT 23.630 8.190 23.860 9.050 ;
        RECT 19.050 7.930 22.250 8.110 ;
        RECT 22.560 8.000 26.230 8.190 ;
        RECT 21.930 7.680 22.110 7.930 ;
        RECT 22.590 7.870 22.820 8.000 ;
        RECT 23.060 7.870 23.290 8.000 ;
        RECT 22.795 7.680 23.085 7.710 ;
        RECT 21.930 7.500 23.085 7.680 ;
        RECT 22.795 7.480 23.085 7.500 ;
        RECT 23.630 7.110 23.860 8.000 ;
        RECT 11.600 6.630 12.450 6.810 ;
        RECT 11.600 6.560 11.830 6.630 ;
        RECT 12.270 6.440 12.450 6.630 ;
        RECT 11.930 6.260 12.450 6.440 ;
        RECT 11.930 5.890 12.110 6.260 ;
        RECT 10.700 5.660 12.260 5.890 ;
        RECT 26.040 5.615 26.230 8.000 ;
        RECT 34.715 5.615 34.905 11.795 ;
        RECT 26.040 5.425 34.905 5.615 ;
        RECT 26.040 2.450 26.230 5.425 ;
        RECT 26.005 2.130 26.265 2.450 ;
        RECT 25.975 0.960 26.295 1.220 ;
        RECT 26.040 0.410 26.230 0.960 ;
        RECT 23.795 0.180 29.865 0.410 ;
      LAYER met2 ;
        RECT 59.425 63.910 59.895 63.930 ;
        RECT 59.400 63.390 62.100 63.910 ;
        RECT 59.425 63.370 59.895 63.390 ;
        RECT 12.080 32.130 12.400 32.390 ;
        RECT 12.110 31.020 12.370 32.130 ;
        RECT 13.380 31.310 13.640 31.340 ;
        RECT 13.380 31.050 14.950 31.310 ;
        RECT 13.380 31.020 13.640 31.050 ;
        RECT 13.820 29.300 14.080 29.620 ;
        RECT 13.870 28.010 14.030 29.300 ;
        RECT 13.790 27.750 14.110 28.010 ;
        RECT 23.650 27.680 23.970 27.940 ;
        RECT 25.670 27.890 25.990 28.150 ;
        RECT 23.695 26.030 23.925 27.680 ;
        RECT 25.740 26.920 25.920 27.890 ;
        RECT 25.700 26.600 25.960 26.920 ;
        RECT 23.650 25.770 23.970 26.030 ;
        RECT 11.250 25.590 11.510 25.670 ;
        RECT 12.410 25.590 12.730 25.640 ;
        RECT 1.130 25.230 1.390 25.550 ;
        RECT 11.250 25.430 12.730 25.590 ;
        RECT 11.250 25.350 11.510 25.430 ;
        RECT 12.410 25.380 12.730 25.430 ;
        RECT 1.150 24.160 1.370 25.230 ;
        RECT 1.130 23.840 1.390 24.160 ;
        RECT 12.330 11.810 12.590 11.880 ;
        RECT 13.250 11.810 13.570 11.850 ;
        RECT 12.330 11.630 13.570 11.810 ;
        RECT 12.330 11.560 12.590 11.630 ;
        RECT 13.250 11.590 13.570 11.630 ;
        RECT 1.870 10.640 2.190 10.900 ;
        RECT 1.935 9.870 2.125 10.640 ;
        RECT 12.200 10.390 12.520 10.650 ;
        RECT 1.900 9.550 2.160 9.870 ;
        RECT 12.270 9.710 12.450 10.390 ;
        RECT 12.230 9.390 12.490 9.710 ;
        RECT 25.975 2.160 26.295 2.420 ;
        RECT 26.040 1.250 26.230 2.160 ;
        RECT 26.005 0.930 26.265 1.250 ;
      LAYER met3 ;
        RECT 57.145 63.910 57.655 63.935 ;
        RECT 57.140 63.390 59.920 63.910 ;
        RECT 57.145 63.365 57.655 63.390 ;
      LAYER met4 ;
        RECT -327.460 427.570 -322.290 427.630 ;
        RECT -321.825 427.570 -292.215 442.115 ;
        RECT -290.225 427.570 -260.615 442.115 ;
        RECT -258.625 427.570 -229.015 442.115 ;
        RECT -227.025 427.570 -197.415 442.115 ;
        RECT -195.425 427.570 -165.815 442.115 ;
        RECT -163.825 427.570 -134.215 442.115 ;
        RECT -132.225 427.570 -102.615 442.115 ;
        RECT -100.625 427.570 -71.015 442.115 ;
        RECT -69.025 427.570 -39.415 442.115 ;
        RECT -37.425 427.570 -7.815 442.115 ;
        RECT -5.825 427.570 23.785 442.115 ;
        RECT 25.775 427.570 55.385 442.115 ;
        RECT -327.460 427.110 56.380 427.570 ;
        RECT -327.460 394.510 -326.940 427.110 ;
        RECT -322.820 427.050 56.380 427.110 ;
        RECT -321.825 412.505 -292.215 427.050 ;
        RECT -290.225 412.505 -260.615 427.050 ;
        RECT -258.625 412.505 -229.015 427.050 ;
        RECT -227.025 412.505 -197.415 427.050 ;
        RECT -195.425 412.505 -165.815 427.050 ;
        RECT -163.825 412.505 -134.215 427.050 ;
        RECT -132.225 412.505 -102.615 427.050 ;
        RECT -100.625 412.505 -71.015 427.050 ;
        RECT -69.025 412.505 -39.415 427.050 ;
        RECT -37.425 412.505 -7.815 427.050 ;
        RECT -5.825 412.505 23.785 427.050 ;
        RECT 25.775 412.505 55.385 427.050 ;
        RECT -321.825 394.510 -292.215 409.055 ;
        RECT -290.225 394.510 -260.615 409.055 ;
        RECT -258.625 394.510 -229.015 409.055 ;
        RECT -227.025 394.510 -197.415 409.055 ;
        RECT -195.425 394.510 -165.815 409.055 ;
        RECT -163.825 394.510 -134.215 409.055 ;
        RECT -132.225 394.510 -102.615 409.055 ;
        RECT -100.625 394.510 -71.015 409.055 ;
        RECT -69.025 394.510 -39.415 409.055 ;
        RECT -37.425 394.510 -7.815 409.055 ;
        RECT -5.825 394.510 23.785 409.055 ;
        RECT 25.775 394.510 55.385 409.055 ;
        RECT -327.460 394.490 56.380 394.510 ;
        RECT -327.460 393.990 59.910 394.490 ;
        RECT -321.825 379.445 -292.215 393.990 ;
        RECT -290.225 379.445 -260.615 393.990 ;
        RECT -258.625 379.445 -229.015 393.990 ;
        RECT -227.025 379.445 -197.415 393.990 ;
        RECT -195.425 379.445 -165.815 393.990 ;
        RECT -163.825 379.445 -134.215 393.990 ;
        RECT -132.225 379.445 -102.615 393.990 ;
        RECT -100.625 379.445 -71.015 393.990 ;
        RECT -69.025 379.445 -39.415 393.990 ;
        RECT -37.425 379.445 -7.815 393.990 ;
        RECT -5.825 379.445 23.785 393.990 ;
        RECT 25.775 379.445 55.385 393.990 ;
        RECT 55.920 393.970 59.910 393.990 ;
        RECT -321.825 361.450 -292.215 375.995 ;
        RECT -290.225 361.450 -260.615 375.995 ;
        RECT -258.625 361.450 -229.015 375.995 ;
        RECT -227.025 361.450 -197.415 375.995 ;
        RECT -195.425 361.450 -165.815 375.995 ;
        RECT -163.825 361.450 -134.215 375.995 ;
        RECT -132.225 361.450 -102.615 375.995 ;
        RECT -100.625 361.450 -71.015 375.995 ;
        RECT -69.025 361.450 -39.415 375.995 ;
        RECT -37.425 361.450 -7.815 375.995 ;
        RECT -5.825 361.450 23.785 375.995 ;
        RECT 25.775 361.450 55.385 375.995 ;
        RECT 59.390 361.450 59.910 393.970 ;
        RECT -322.820 361.400 59.910 361.450 ;
        RECT -326.020 360.930 59.910 361.400 ;
        RECT -326.020 360.880 -322.250 360.930 ;
        RECT -326.020 328.390 -325.500 360.880 ;
        RECT -321.825 346.385 -292.215 360.930 ;
        RECT -290.225 346.385 -260.615 360.930 ;
        RECT -258.625 346.385 -229.015 360.930 ;
        RECT -227.025 346.385 -197.415 360.930 ;
        RECT -195.425 346.385 -165.815 360.930 ;
        RECT -163.825 346.385 -134.215 360.930 ;
        RECT -132.225 346.385 -102.615 360.930 ;
        RECT -100.625 346.385 -71.015 360.930 ;
        RECT -69.025 346.385 -39.415 360.930 ;
        RECT -37.425 346.385 -7.815 360.930 ;
        RECT -5.825 346.385 23.785 360.930 ;
        RECT 25.775 346.385 55.385 360.930 ;
        RECT -321.825 328.390 -292.215 342.935 ;
        RECT -290.225 328.390 -260.615 342.935 ;
        RECT -258.625 328.390 -229.015 342.935 ;
        RECT -227.025 328.390 -197.415 342.935 ;
        RECT -195.425 328.390 -165.815 342.935 ;
        RECT -163.825 328.390 -134.215 342.935 ;
        RECT -132.225 328.390 -102.615 342.935 ;
        RECT -100.625 328.390 -71.015 342.935 ;
        RECT -69.025 328.390 -39.415 342.935 ;
        RECT -37.425 328.390 -7.815 342.935 ;
        RECT -5.825 328.390 23.785 342.935 ;
        RECT 25.775 328.390 55.385 342.935 ;
        RECT -326.020 328.350 56.380 328.390 ;
        RECT -326.020 327.870 61.220 328.350 ;
        RECT -321.825 313.325 -292.215 327.870 ;
        RECT -290.225 313.325 -260.615 327.870 ;
        RECT -258.625 313.325 -229.015 327.870 ;
        RECT -227.025 313.325 -197.415 327.870 ;
        RECT -195.425 313.325 -165.815 327.870 ;
        RECT -163.825 313.325 -134.215 327.870 ;
        RECT -132.225 313.325 -102.615 327.870 ;
        RECT -100.625 313.325 -71.015 327.870 ;
        RECT -69.025 313.325 -39.415 327.870 ;
        RECT -37.425 313.325 -7.815 327.870 ;
        RECT -5.825 313.325 23.785 327.870 ;
        RECT 25.775 313.325 55.385 327.870 ;
        RECT 56.030 327.830 61.220 327.870 ;
        RECT -325.290 295.330 -322.250 295.420 ;
        RECT -321.825 295.330 -292.215 309.875 ;
        RECT -290.225 295.330 -260.615 309.875 ;
        RECT -258.625 295.330 -229.015 309.875 ;
        RECT -227.025 295.330 -197.415 309.875 ;
        RECT -195.425 295.330 -165.815 309.875 ;
        RECT -163.825 295.330 -134.215 309.875 ;
        RECT -132.225 295.330 -102.615 309.875 ;
        RECT -100.625 295.330 -71.015 309.875 ;
        RECT -69.025 295.330 -39.415 309.875 ;
        RECT -37.425 295.330 -7.815 309.875 ;
        RECT -5.825 295.330 23.785 309.875 ;
        RECT 25.775 295.330 55.385 309.875 ;
        RECT 60.700 295.330 61.220 327.830 ;
        RECT -325.290 294.900 61.220 295.330 ;
        RECT -325.290 262.270 -324.770 294.900 ;
        RECT -322.820 294.810 61.220 294.900 ;
        RECT -321.825 280.265 -292.215 294.810 ;
        RECT -290.225 280.265 -260.615 294.810 ;
        RECT -258.625 280.265 -229.015 294.810 ;
        RECT -227.025 280.265 -197.415 294.810 ;
        RECT -195.425 280.265 -165.815 294.810 ;
        RECT -163.825 280.265 -134.215 294.810 ;
        RECT -132.225 280.265 -102.615 294.810 ;
        RECT -100.625 280.265 -71.015 294.810 ;
        RECT -69.025 280.265 -39.415 294.810 ;
        RECT -37.425 280.265 -7.815 294.810 ;
        RECT -5.825 280.265 23.785 294.810 ;
        RECT 25.775 280.265 55.385 294.810 ;
        RECT -321.825 262.270 -292.215 276.815 ;
        RECT -290.225 262.270 -260.615 276.815 ;
        RECT -258.625 262.270 -229.015 276.815 ;
        RECT -227.025 262.270 -197.415 276.815 ;
        RECT -195.425 262.270 -165.815 276.815 ;
        RECT -163.825 262.270 -134.215 276.815 ;
        RECT -132.225 262.270 -102.615 276.815 ;
        RECT -100.625 262.270 -71.015 276.815 ;
        RECT -69.025 262.270 -39.415 276.815 ;
        RECT -37.425 262.270 -7.815 276.815 ;
        RECT -5.825 262.270 23.785 276.815 ;
        RECT 25.775 262.270 55.385 276.815 ;
        RECT 55.870 262.270 60.480 262.310 ;
        RECT -325.290 261.790 60.480 262.270 ;
        RECT -325.290 261.750 56.380 261.790 ;
        RECT -321.825 247.205 -292.215 261.750 ;
        RECT -290.225 247.205 -260.615 261.750 ;
        RECT -258.625 247.205 -229.015 261.750 ;
        RECT -227.025 247.205 -197.415 261.750 ;
        RECT -195.425 247.205 -165.815 261.750 ;
        RECT -163.825 247.205 -134.215 261.750 ;
        RECT -132.225 247.205 -102.615 261.750 ;
        RECT -100.625 247.205 -71.015 261.750 ;
        RECT -69.025 247.205 -39.415 261.750 ;
        RECT -37.425 247.205 -7.815 261.750 ;
        RECT -5.825 247.205 23.785 261.750 ;
        RECT 25.775 247.205 55.385 261.750 ;
        RECT -321.825 229.210 -292.215 243.755 ;
        RECT -290.225 229.210 -260.615 243.755 ;
        RECT -258.625 229.210 -229.015 243.755 ;
        RECT -227.025 229.210 -197.415 243.755 ;
        RECT -195.425 229.210 -165.815 243.755 ;
        RECT -163.825 229.210 -134.215 243.755 ;
        RECT -132.225 229.210 -102.615 243.755 ;
        RECT -100.625 229.210 -71.015 243.755 ;
        RECT -69.025 229.210 -39.415 243.755 ;
        RECT -37.425 229.210 -7.815 243.755 ;
        RECT -5.825 229.210 23.785 243.755 ;
        RECT 25.775 229.210 55.385 243.755 ;
        RECT 59.960 229.210 60.480 261.790 ;
        RECT -327.630 228.690 60.480 229.210 ;
        RECT -327.630 196.150 -327.110 228.690 ;
        RECT -321.825 214.145 -292.215 228.690 ;
        RECT -290.225 214.145 -260.615 228.690 ;
        RECT -258.625 214.145 -229.015 228.690 ;
        RECT -227.025 214.145 -197.415 228.690 ;
        RECT -195.425 214.145 -165.815 228.690 ;
        RECT -163.825 214.145 -134.215 228.690 ;
        RECT -132.225 214.145 -102.615 228.690 ;
        RECT -100.625 214.145 -71.015 228.690 ;
        RECT -69.025 214.145 -39.415 228.690 ;
        RECT -37.425 214.145 -7.815 228.690 ;
        RECT -5.825 214.145 23.785 228.690 ;
        RECT 25.775 214.145 55.385 228.690 ;
        RECT -321.825 196.150 -292.215 210.695 ;
        RECT -290.225 196.150 -260.615 210.695 ;
        RECT -258.625 196.150 -229.015 210.695 ;
        RECT -227.025 196.150 -197.415 210.695 ;
        RECT -195.425 196.150 -165.815 210.695 ;
        RECT -163.825 196.150 -134.215 210.695 ;
        RECT -132.225 196.150 -102.615 210.695 ;
        RECT -100.625 196.150 -71.015 210.695 ;
        RECT -69.025 196.150 -39.415 210.695 ;
        RECT -37.425 196.150 -7.815 210.695 ;
        RECT -5.825 196.150 23.785 210.695 ;
        RECT 25.775 196.150 55.385 210.695 ;
        RECT 55.910 196.150 58.930 196.160 ;
        RECT -327.630 195.640 58.930 196.150 ;
        RECT -327.630 195.630 56.380 195.640 ;
        RECT -321.825 181.085 -292.215 195.630 ;
        RECT -290.225 181.085 -260.615 195.630 ;
        RECT -258.625 181.085 -229.015 195.630 ;
        RECT -227.025 181.085 -197.415 195.630 ;
        RECT -195.425 181.085 -165.815 195.630 ;
        RECT -163.825 181.085 -134.215 195.630 ;
        RECT -132.225 181.085 -102.615 195.630 ;
        RECT -100.625 181.085 -71.015 195.630 ;
        RECT -69.025 181.085 -39.415 195.630 ;
        RECT -37.425 181.085 -7.815 195.630 ;
        RECT -5.825 181.085 23.785 195.630 ;
        RECT 25.775 181.085 55.385 195.630 ;
        RECT -321.825 163.090 -292.215 177.635 ;
        RECT -290.225 163.090 -260.615 177.635 ;
        RECT -258.625 163.090 -229.015 177.635 ;
        RECT -227.025 163.090 -197.415 177.635 ;
        RECT -195.425 163.090 -165.815 177.635 ;
        RECT -163.825 163.090 -134.215 177.635 ;
        RECT -132.225 163.090 -102.615 177.635 ;
        RECT -100.625 163.090 -71.015 177.635 ;
        RECT -69.025 163.090 -39.415 177.635 ;
        RECT -37.425 163.090 -7.815 177.635 ;
        RECT -5.825 163.090 23.785 177.635 ;
        RECT 25.775 163.090 55.385 177.635 ;
        RECT 58.410 163.090 58.930 195.640 ;
        RECT -322.820 163.030 58.930 163.090 ;
        RECT -326.150 162.570 58.930 163.030 ;
        RECT -326.150 162.510 -322.270 162.570 ;
        RECT -326.150 130.030 -325.630 162.510 ;
        RECT -321.825 148.025 -292.215 162.570 ;
        RECT -290.225 148.025 -260.615 162.570 ;
        RECT -258.625 148.025 -229.015 162.570 ;
        RECT -227.025 148.025 -197.415 162.570 ;
        RECT -195.425 148.025 -165.815 162.570 ;
        RECT -163.825 148.025 -134.215 162.570 ;
        RECT -132.225 148.025 -102.615 162.570 ;
        RECT -100.625 148.025 -71.015 162.570 ;
        RECT -69.025 148.025 -39.415 162.570 ;
        RECT -37.425 148.025 -7.815 162.570 ;
        RECT -5.825 148.025 23.785 162.570 ;
        RECT 25.775 148.025 55.385 162.570 ;
        RECT -321.825 130.030 -292.215 144.575 ;
        RECT -290.225 130.030 -260.615 144.575 ;
        RECT -258.625 130.030 -229.015 144.575 ;
        RECT -227.025 130.030 -197.415 144.575 ;
        RECT -195.425 130.030 -165.815 144.575 ;
        RECT -163.825 130.030 -134.215 144.575 ;
        RECT -132.225 130.030 -102.615 144.575 ;
        RECT -100.625 130.030 -71.015 144.575 ;
        RECT -69.025 130.030 -39.415 144.575 ;
        RECT -37.425 130.030 -7.815 144.575 ;
        RECT -5.825 130.030 23.785 144.575 ;
        RECT 25.775 130.030 55.385 144.575 ;
        RECT -326.150 129.960 56.380 130.030 ;
        RECT -326.150 129.510 59.930 129.960 ;
        RECT -321.825 114.965 -292.215 129.510 ;
        RECT -290.225 114.965 -260.615 129.510 ;
        RECT -258.625 114.965 -229.015 129.510 ;
        RECT -227.025 114.965 -197.415 129.510 ;
        RECT -195.425 114.965 -165.815 129.510 ;
        RECT -163.825 114.965 -134.215 129.510 ;
        RECT -132.225 114.965 -102.615 129.510 ;
        RECT -100.625 114.965 -71.015 129.510 ;
        RECT -69.025 114.965 -39.415 129.510 ;
        RECT -37.425 114.965 -7.815 129.510 ;
        RECT -5.825 114.965 23.785 129.510 ;
        RECT 25.775 114.965 55.385 129.510 ;
        RECT 56.030 129.440 59.930 129.510 ;
        RECT -321.825 96.970 -292.215 111.515 ;
        RECT -290.225 96.970 -260.615 111.515 ;
        RECT -258.625 96.970 -229.015 111.515 ;
        RECT -227.025 96.970 -197.415 111.515 ;
        RECT -195.425 96.970 -165.815 111.515 ;
        RECT -163.825 96.970 -134.215 111.515 ;
        RECT -132.225 96.970 -102.615 111.515 ;
        RECT -100.625 96.970 -71.015 111.515 ;
        RECT -69.025 96.970 -39.415 111.515 ;
        RECT -37.425 96.970 -7.815 111.515 ;
        RECT -5.825 96.970 23.785 111.515 ;
        RECT 25.775 96.970 55.385 111.515 ;
        RECT 59.410 96.970 59.930 129.440 ;
        RECT -322.820 96.820 59.930 96.970 ;
        RECT -326.940 96.450 59.930 96.820 ;
        RECT -326.940 96.300 -322.350 96.450 ;
        RECT -326.940 63.910 -326.420 96.300 ;
        RECT -321.825 81.905 -292.215 96.450 ;
        RECT -290.225 81.905 -260.615 96.450 ;
        RECT -258.625 81.905 -229.015 96.450 ;
        RECT -227.025 81.905 -197.415 96.450 ;
        RECT -195.425 81.905 -165.815 96.450 ;
        RECT -163.825 81.905 -134.215 96.450 ;
        RECT -132.225 81.905 -102.615 96.450 ;
        RECT -100.625 81.905 -71.015 96.450 ;
        RECT -69.025 81.905 -39.415 96.450 ;
        RECT -37.425 81.905 -7.815 96.450 ;
        RECT -5.825 81.905 23.785 96.450 ;
        RECT 25.775 81.905 55.385 96.450 ;
        RECT -321.825 63.910 -292.215 78.455 ;
        RECT -290.225 63.910 -260.615 78.455 ;
        RECT -258.625 63.910 -229.015 78.455 ;
        RECT -227.025 63.910 -197.415 78.455 ;
        RECT -195.425 63.910 -165.815 78.455 ;
        RECT -163.825 63.910 -134.215 78.455 ;
        RECT -132.225 63.910 -102.615 78.455 ;
        RECT -100.625 63.910 -71.015 78.455 ;
        RECT -69.025 63.910 -39.415 78.455 ;
        RECT -37.425 63.910 -7.815 78.455 ;
        RECT -5.825 63.910 23.785 78.455 ;
        RECT 25.775 63.910 55.385 78.455 ;
        RECT -326.940 63.390 57.660 63.910 ;
        RECT -321.825 48.845 -292.215 63.390 ;
        RECT -290.225 48.845 -260.615 63.390 ;
        RECT -258.625 48.845 -229.015 63.390 ;
        RECT -227.025 48.845 -197.415 63.390 ;
        RECT -195.425 48.845 -165.815 63.390 ;
        RECT -163.825 48.845 -134.215 63.390 ;
        RECT -132.225 48.845 -102.615 63.390 ;
        RECT -100.625 48.845 -71.015 63.390 ;
        RECT -69.025 48.845 -39.415 63.390 ;
        RECT -37.425 48.845 -7.815 63.390 ;
        RECT -5.825 48.845 23.785 63.390 ;
        RECT 25.775 48.845 55.385 63.390 ;
  END
END cp
END LIBRARY

