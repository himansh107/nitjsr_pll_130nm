VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__pfet_01v8_X4438S
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__pfet_01v8_X4438S ;
  ORIGIN 0.805 1.190 ;
  SIZE 1.610 BY 2.380 ;
  OBS
      LAYER nwell ;
        RECT -1.070 -1.455 1.070 1.455 ;
      LAYER li1 ;
        RECT -0.890 1.105 0.890 1.275 ;
        RECT -0.890 -1.105 -0.720 1.105 ;
        RECT -0.165 0.595 0.165 0.765 ;
        RECT -0.320 -0.380 -0.150 0.380 ;
        RECT 0.150 -0.380 0.320 0.380 ;
        RECT -0.165 -0.765 0.165 -0.595 ;
        RECT 0.720 -1.105 0.890 1.105 ;
        RECT -0.890 -1.275 0.890 -1.105 ;
      LAYER met1 ;
        RECT -0.145 0.565 0.145 0.795 ;
        RECT -0.350 -0.360 -0.120 0.360 ;
        RECT 0.120 -0.360 0.350 0.360 ;
        RECT -0.145 -0.795 0.145 -0.565 ;
  END
END sky130_fd_pr__pfet_01v8_X4438S
MACRO sky130_fd_pr__nfet_01v8_4BNSKG
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__nfet_01v8_4BNSKG ;
  ORIGIN 0.805 0.995 ;
  SIZE 1.610 BY 1.990 ;
  OBS
      LAYER pwell ;
        RECT -1.070 -1.260 1.070 1.260 ;
      LAYER li1 ;
        RECT -0.890 0.910 0.890 1.080 ;
        RECT -0.890 -0.910 -0.720 0.910 ;
        RECT -0.165 0.400 0.165 0.570 ;
        RECT -0.320 -0.230 -0.150 0.230 ;
        RECT 0.150 -0.230 0.320 0.230 ;
        RECT -0.165 -0.570 0.165 -0.400 ;
        RECT 0.720 -0.910 0.890 0.910 ;
        RECT -0.890 -1.080 0.890 -0.910 ;
      LAYER met1 ;
        RECT -0.145 0.370 0.145 0.600 ;
        RECT -0.350 -0.210 -0.120 0.210 ;
        RECT 0.120 -0.210 0.350 0.210 ;
        RECT -0.145 -0.600 0.145 -0.370 ;
  END
END sky130_fd_pr__nfet_01v8_4BNSKG
MACRO sky130_fd_pr__nfet_01v8_6FB46G
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__nfet_01v8_6FB46G ;
  ORIGIN 0.805 0.995 ;
  SIZE 1.610 BY 1.990 ;
  OBS
      LAYER pwell ;
        RECT -1.070 -1.260 1.070 1.260 ;
      LAYER li1 ;
        RECT -0.890 0.910 0.890 1.080 ;
        RECT -0.890 -0.910 -0.720 0.910 ;
        RECT -0.165 0.400 0.165 0.570 ;
        RECT -0.320 -0.230 -0.150 0.230 ;
        RECT 0.150 -0.230 0.320 0.230 ;
        RECT -0.165 -0.570 0.165 -0.400 ;
        RECT 0.720 -0.910 0.890 0.910 ;
        RECT -0.890 -1.080 0.890 -0.910 ;
      LAYER met1 ;
        RECT -0.145 0.370 0.145 0.600 ;
        RECT -0.350 -0.210 -0.120 0.210 ;
        RECT 0.120 -0.210 0.350 0.210 ;
        RECT -0.145 -0.600 0.145 -0.370 ;
        RECT -0.780 -1.110 0.780 -0.880 ;
  END
END sky130_fd_pr__nfet_01v8_6FB46G
MACRO cs_inv
  CLASS BLOCK ;
  FOREIGN cs_inv ;
  ORIGIN -1.465 10.190 ;
  SIZE 6.890 BY 13.070 ;
  PIN Vp
    ANTENNAGATEAREA 0.129600 ;
    PORT
      LAYER li1 ;
        RECT 5.230 0.770 5.560 0.940 ;
        RECT 5.230 -0.590 5.560 -0.420 ;
      LAYER met1 ;
        RECT 5.250 0.920 5.540 0.970 ;
        RECT 3.765 0.770 5.540 0.920 ;
        RECT 2.105 0.340 3.105 0.700 ;
        RECT 3.775 0.340 3.965 0.770 ;
        RECT 5.250 0.740 5.540 0.770 ;
        RECT 2.105 0.070 3.965 0.340 ;
        RECT 2.105 -0.300 3.105 0.070 ;
        RECT 3.775 -0.430 3.965 0.070 ;
        RECT 5.250 -0.430 5.540 -0.390 ;
        RECT 3.775 -0.580 5.565 -0.430 ;
        RECT 5.250 -0.620 5.540 -0.580 ;
    END
  END Vp
  PIN out
    ANTENNADIFFAREA 0.330600 ;
    PORT
      LAYER li1 ;
        RECT 5.545 -3.025 5.715 -2.265 ;
        RECT 5.085 -5.830 5.255 -5.370 ;
      LAYER met1 ;
        RECT 5.515 -2.790 5.745 -2.285 ;
        RECT 6.515 -2.790 6.695 -2.785 ;
        RECT 5.515 -2.960 6.705 -2.790 ;
        RECT 5.515 -3.005 5.745 -2.960 ;
        RECT 6.515 -3.750 6.695 -2.960 ;
        RECT 7.355 -3.750 8.355 -3.350 ;
        RECT 6.505 -3.970 8.355 -3.750 ;
        RECT 4.295 -4.470 4.615 -4.430 ;
        RECT 6.515 -4.470 6.695 -3.970 ;
        RECT 7.355 -4.350 8.355 -3.970 ;
        RECT 4.295 -4.650 6.695 -4.470 ;
        RECT 4.295 -4.690 4.615 -4.650 ;
        RECT 6.515 -4.670 6.695 -4.650 ;
        RECT 4.325 -5.460 4.585 -5.390 ;
        RECT 5.055 -5.460 5.285 -5.390 ;
        RECT 4.325 -5.640 5.285 -5.460 ;
        RECT 4.325 -5.710 4.585 -5.640 ;
        RECT 4.905 -5.650 5.285 -5.640 ;
      