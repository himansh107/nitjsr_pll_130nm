magic
tech sky130A
magscale 1 2
timestamp 1713377695
<< error_p >>
rect -29 331 29 337
rect -29 297 -17 331
rect -29 291 29 297
rect -29 -297 29 -291
rect -29 -331 -17 -297
rect -29 -337 29 -331
<< nwell >>
rect -211 -469 211 469
<< pmos >>
rect -15 -250 15 250
<< pdiff >>
rect -73 238 -15 250
rect -73 -238 -61 238
rect -27 -238 -15 238
rect -73 -250 -15 -238
rect 15 238 73 250
rect 15 -238 27 238
rect 61 -238 73 238
rect 15 -250 73 -238
<< pdiffc >>
rect -61 -238 -27 238
rect 27 -238 61 238
<< nsubdiff >>
rect -175 399 -79 433
rect 79 399 175 433
rect -175 337 -141 399
rect 141 337 175 399
rect -175 -399 -141 -337
rect 141 -399 175 -337
rect -175 -433 -79 -399
rect 79 -433 175 -399
<< nsubdiffcont >>
rect -79 399 79 433
rect -175 -337 -141 337
rect 141 -337 175 337
rect -79 -433 79 -399
<< poly >>
rect -33 331 33 347
rect -33 297 -17 331
rect 17 297 33 331
rect -33 281 33 297
rect -15 250 15 281
rect -15 -281 15 -250
rect -33 -297 33 -281
rect -33 -331 -17 -297
rect 17 -331 33 -297
rect -33 -347 33 -331
<< polycont >>
rect -17 297 17 331
rect -17 -331 17 -297
<< locali >>
rect -175 399 -79 433
rect 79 399 175 433
rect -175 337 -141 399
rect 141 337 175 399
rect -33 297 -17 331
rect 17 297 33 331
rect -61 238 -27 254
rect -61 -254 -27 -238
rect 27 238 61 254
rect 27 -254 61 -238
rect -33 -331 -17 -297
rect 17 -331 33 -297
rect -175 -399 -141 -337
rect 141 -399 175 -337
rect -175 -433 -79 -399
rect 79 -433 175 -399
<< viali >>
rect -17 297 17 331
rect -61 -238 -27 238
rect 27 -238 61 238
rect -17 -331 17 -297
<< metal1 >>
rect -29 331 29 337
rect -29 297 -17 331
rect 17 297 29 331
rect -29 291 29 297
rect -67 238 -21 250
rect -67 -238 -61 238
rect -27 -238 -21 238
rect -67 -250 -21 -238
rect 21 238 67 250
rect 21 -238 27 238
rect 61 -238 67 238
rect 21 -250 67 -238
rect -29 -297 29 -291
rect -29 -331 -17 -297
rect 17 -331 29 -297
rect -29 -337 29 -331
<< properties >>
string FIXED_BBOX -158 -416 158 416
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
