magic
tech sky130A
magscale 1 2
timestamp 1714283992
<< error_p >>
rect -29 4581 29 4587
rect -29 4547 -17 4581
rect -29 4541 29 4547
rect -29 -4547 29 -4541
rect -29 -4581 -17 -4547
rect -29 -4587 29 -4581
<< nwell >>
rect -214 -4719 214 4719
<< pmos >>
rect -18 -4500 18 4500
<< pdiff >>
rect -76 4488 -18 4500
rect -76 -4488 -64 4488
rect -30 -4488 -18 4488
rect -76 -4500 -18 -4488
rect 18 4488 76 4500
rect 18 -4488 30 4488
rect 64 -4488 76 4488
rect 18 -4500 76 -4488
<< pdiffc >>
rect -64 -4488 -30 4488
rect 30 -4488 64 4488
<< nsubdiff >>
rect -178 4649 -82 4683
rect 82 4649 178 4683
rect -178 4587 -144 4649
rect 144 4587 178 4649
rect -178 -4649 -144 -4587
rect 144 -4649 178 -4587
rect -178 -4683 -82 -4649
rect 82 -4683 178 -4649
<< nsubdiffcont >>
rect -82 4649 82 4683
rect -178 -4587 -144 4587
rect 144 -4587 178 4587
rect -82 -4683 82 -4649
<< poly >>
rect -33 4581 33 4597
rect -33 4547 -17 4581
rect 17 4547 33 4581
rect -33 4531 33 4547
rect -18 4500 18 4531
rect -18 -4531 18 -4500
rect -33 -4547 33 -4531
rect -33 -4581 -17 -4547
rect 17 -4581 33 -4547
rect -33 -4597 33 -4581
<< polycont >>
rect -17 4547 17 4581
rect -17 -4581 17 -4547
<< locali >>
rect -178 4587 -144 4683
rect 144 4587 178 4683
rect -33 4547 -17 4581
rect 17 4547 33 4581
rect -64 4488 -30 4504
rect -64 -4504 -30 -4488
rect 30 4488 64 4504
rect 30 -4504 64 -4488
rect -33 -4581 -17 -4547
rect 17 -4581 33 -4547
rect -178 -4649 -144 -4587
rect 144 -4649 178 -4587
rect -178 -4683 -82 -4649
rect 82 -4683 178 -4649
<< viali >>
rect -144 4649 -82 4683
rect -82 4649 82 4683
rect 82 4649 144 4683
rect -17 4547 17 4581
rect -64 881 -30 4471
rect 30 -4471 64 -881
rect -17 -4581 17 -4547
<< metal1 >>
rect -156 4683 156 4689
rect -156 4649 -144 4683
rect 144 4649 156 4683
rect -156 4643 156 4649
rect -29 4581 29 4587
rect -29 4547 -17 4581
rect 17 4547 29 4581
rect -29 4541 29 4547
rect -70 4471 -24 4483
rect -70 881 -64 4471
rect -30 881 -24 4471
rect -70 869 -24 881
rect 24 -881 70 -869
rect 24 -4471 30 -881
rect 64 -4471 70 -881
rect 24 -4483 70 -4471
rect -29 -4547 29 -4541
rect -29 -4581 -17 -4547
rect 17 -4581 29 -4547
rect -29 -4587 29 -4581
<< properties >>
string FIXED_BBOX -161 -4666 161 4666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 45.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
