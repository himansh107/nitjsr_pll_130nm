magic
tech sky130A
magscale 1 2
timestamp 1713777229
<< pwell >>
rect 13588 -3878 13790 -3828
<< viali >>
rect 13618 -2768 13786 -2730
rect 13588 -3878 13790 -3828
<< metal1 >>
rect 2594 -1788 2648 -1786
rect 4114 -1788 4168 -1778
rect 5644 -1788 5698 -1786
rect 7212 -1788 7266 -1778
rect 8796 -1788 8850 -1786
rect 10330 -1788 10384 -1784
rect 2352 -1842 11844 -1788
rect 1852 -2091 1898 -2082
rect 2240 -2091 2246 -2088
rect 1852 -2137 2246 -2091
rect 1852 -2218 1898 -2137
rect 2240 -2140 2246 -2137
rect 2298 -2140 2304 -2088
rect 1766 -2536 1966 -2218
rect 1816 -2662 1864 -2536
rect 1382 -2702 1864 -2662
rect 1098 -2766 1478 -2764
rect 1096 -2816 1478 -2766
rect 1096 -3250 1142 -2816
rect 1816 -2890 1864 -2702
rect 1384 -2938 1864 -2890
rect 1472 -3180 1706 -3154
rect 2352 -3179 2406 -1842
rect 2594 -2668 2648 -1842
rect 2726 -2088 2778 -2082
rect 3952 -2091 3958 -2088
rect 2778 -2137 3958 -2091
rect 3952 -2140 3958 -2137
rect 4010 -2140 4016 -2088
rect 2726 -2146 2778 -2140
rect 4114 -2660 4168 -1842
rect 4264 -2088 4316 -2082
rect 5516 -2091 5522 -2088
rect 4316 -2137 5522 -2091
rect 5516 -2140 5522 -2137
rect 5574 -2140 5580 -2088
rect 4264 -2146 4316 -2140
rect 5644 -2668 5698 -1842
rect 5752 -2088 5804 -2082
rect 7112 -2088 7164 -2082
rect 5804 -2137 7112 -2091
rect 5752 -2146 5804 -2140
rect 7112 -2146 7164 -2140
rect 7212 -2660 7266 -1842
rect 7336 -2088 7388 -2082
rect 8634 -2091 8640 -2088
rect 7388 -2137 8640 -2091
rect 8634 -2140 8640 -2137
rect 8692 -2140 8698 -2088
rect 7336 -2146 7388 -2140
rect 8796 -2668 8850 -1842
rect 8910 -2088 8962 -2082
rect 10220 -2091 10226 -2088
rect 8962 -2137 10226 -2091
rect 10220 -2140 10226 -2137
rect 10278 -2140 10284 -2088
rect 8910 -2146 8962 -2140
rect 10330 -2666 10384 -1842
rect 10462 -2088 10514 -2082
rect 11666 -2091 11672 -2088
rect 10514 -2137 11672 -2091
rect 11666 -2140 11672 -2137
rect 11724 -2140 11730 -2088
rect 10462 -2146 10514 -2140
rect 11790 -2567 11844 -1842
rect 11882 -2088 11934 -2082
rect 11934 -2137 12425 -2091
rect 11882 -2146 11934 -2140
rect 12468 -2142 13703 -2092
rect 13653 -2480 13703 -2142
rect 13598 -2626 13798 -2480
rect 13422 -2726 13428 -2674
rect 13480 -2682 13486 -2674
rect 13526 -2682 13872 -2626
rect 13480 -2718 13872 -2682
rect 13480 -2726 13486 -2718
rect 13526 -2730 13872 -2718
rect 13526 -2768 13618 -2730
rect 13786 -2768 13872 -2730
rect 13526 -2780 13872 -2768
rect 13302 -2886 13730 -2848
rect 13304 -2968 13340 -2886
rect 13184 -3018 13340 -2968
rect 1798 -3180 2406 -3179
rect 1472 -3194 2406 -3180
rect 1658 -3233 2406 -3194
rect 1096 -3302 1478 -3250
rect 1096 -3479 1142 -3302
rect 1658 -3479 1700 -3233
rect 1096 -3525 1700 -3479
rect 1244 -3638 1250 -3586
rect 1302 -3591 1308 -3586
rect 1658 -3591 1700 -3525
rect 1302 -3633 1700 -3591
rect 1302 -3638 1308 -3633
rect 2467 -3677 2521 -3417
rect 3688 -3436 4104 -3364
rect 5218 -3408 5634 -3336
rect 6690 -3408 7106 -3336
rect 13186 -3344 13220 -3018
rect 13304 -3116 13340 -3018
rect 13428 -2970 13480 -2964
rect 13480 -3014 13662 -2978
rect 13726 -3018 13962 -2980
rect 13428 -3028 13480 -3022
rect 13304 -3154 13732 -3116
rect 8296 -3416 8712 -3344
rect 9884 -3416 10300 -3344
rect 11362 -3426 11778 -3354
rect 12934 -3398 13220 -3344
rect 13923 -3238 13961 -3018
rect 14054 -3238 14254 -3140
rect 13923 -3290 14254 -3238
rect 2085 -3731 2521 -3677
rect 442 -3864 642 -3780
rect 1106 -3782 1474 -3736
rect 1110 -3845 1150 -3782
rect 1003 -3864 1150 -3845
rect 442 -3899 1150 -3864
rect 1244 -3880 1250 -3828
rect 1302 -3833 1308 -3828
rect 1302 -3875 1407 -3833
rect 1302 -3880 1308 -3875
rect 1468 -3890 1716 -3846
rect 442 -3918 1057 -3899
rect 442 -3980 642 -3918
rect 1003 -4788 1057 -3918
rect 1110 -3930 1150 -3899
rect 1108 -3976 1476 -3930
rect 1280 -4108 1602 -4050
rect 1672 -4108 1716 -3890
rect 1280 -4152 1716 -4108
rect 1280 -4224 1602 -4152
rect 1336 -4350 1536 -4224
rect 1452 -4546 1500 -4350
rect 1970 -4546 1976 -4544
rect 1452 -4594 1976 -4546
rect 1970 -4596 1976 -4594
rect 2028 -4596 2034 -4544
rect 1785 -4788 1839 -4782
rect 1003 -4842 1785 -4788
rect 1785 -4848 1839 -4842
rect 2085 -4939 2139 -3731
rect 2220 -4544 2272 -4538
rect 2542 -4546 2548 -4544
rect 2272 -4594 2548 -4546
rect 2542 -4596 2548 -4594
rect 2600 -4596 2606 -4544
rect 2220 -4602 2272 -4596
rect 2650 -4788 2704 -4120
rect 2774 -4544 2826 -4538
rect 4056 -4546 4062 -4544
rect 2826 -4594 4062 -4546
rect 4056 -4596 4062 -4594
rect 4114 -4596 4120 -4544
rect 2774 -4602 2826 -4596
rect 4170 -4788 4224 -4110
rect 4294 -4544 4346 -4538
rect 5578 -4546 5584 -4544
rect 4346 -4594 5584 -4546
rect 5578 -4596 5584 -4594
rect 5636 -4596 5642 -4544
rect 4294 -4602 4346 -4596
rect 5706 -4788 5760 -4108
rect 5854 -4544 5906 -4538
rect 7154 -4546 7160 -4544
rect 5906 -4594 7160 -4546
rect 7154 -4596 7160 -4594
rect 7212 -4596 7218 -4544
rect 5854 -4602 5906 -4596
rect 7282 -4788 7336 -4114
rect 7450 -4544 7502 -4538
rect 8728 -4546 8734 -4544
rect 7502 -4594 8734 -4546
rect 8728 -4596 8734 -4594
rect 8786 -4596 8792 -4544
rect 7450 -4602 7502 -4596
rect 8872 -4788 8926 -4116
rect 8982 -4544 9034 -4538
rect 10316 -4546 10322 -4544
rect 9034 -4594 10322 -4546
rect 10316 -4596 10322 -4594
rect 10374 -4596 10380 -4544
rect 8982 -4602 9034 -4596
rect 10416 -4788 10470 -4116
rect 10556 -4544 10608 -4538
rect 11766 -4546 11772 -4544
rect 10608 -4594 11772 -4546
rect 11766 -4596 11772 -4594
rect 11824 -4596 11830 -4544
rect 10556 -4602 10608 -4596
rect 11900 -4788 11954 -4197
rect 12010 -4544 12062 -4538
rect 12890 -4546 12896 -4544
rect 12062 -4594 12896 -4546
rect 12890 -4596 12896 -4594
rect 12948 -4596 12954 -4544
rect 12010 -4602 12062 -4596
rect 2311 -4842 2317 -4788
rect 2371 -4842 11954 -4788
rect 2650 -4848 2704 -4842
rect 8872 -4844 8926 -4842
rect 10416 -4844 10470 -4842
rect 13025 -4939 13079 -3398
rect 13186 -3598 13220 -3398
rect 13462 -3436 13468 -3384
rect 13520 -3391 13526 -3384
rect 13923 -3391 13961 -3290
rect 14054 -3340 14254 -3290
rect 13520 -3429 13961 -3391
rect 13520 -3436 13526 -3429
rect 13296 -3526 13724 -3524
rect 13290 -3562 13724 -3526
rect 13290 -3598 13332 -3562
rect 13186 -3634 13332 -3598
rect 13188 -3638 13332 -3634
rect 13290 -3720 13332 -3638
rect 13468 -3624 13520 -3618
rect 13520 -3669 13659 -3631
rect 13714 -3666 13928 -3632
rect 13468 -3682 13520 -3676
rect 13290 -3758 13720 -3720
rect 13502 -3828 13858 -3822
rect 13502 -3878 13588 -3828
rect 13790 -3878 13858 -3828
rect 13502 -3893 13858 -3878
rect 13891 -3893 13925 -3666
rect 13502 -3927 13925 -3893
rect 13502 -3986 13858 -3927
rect 13592 -4136 13792 -3986
rect 13314 -4544 13366 -4538
rect 13684 -4546 13732 -4136
rect 13366 -4594 13734 -4546
rect 13314 -4602 13366 -4596
rect 2085 -4993 13079 -4939
<< via1 >>
rect 2246 -2140 2298 -2088
rect 2726 -2140 2778 -2088
rect 3958 -2140 4010 -2088
rect 4264 -2140 4316 -2088
rect 5522 -2140 5574 -2088
rect 5752 -2140 5804 -2088
rect 7112 -2140 7164 -2088
rect 7336 -2140 7388 -2088
rect 8640 -2140 8692 -2088
rect 8910 -2140 8962 -2088
rect 10226 -2140 10278 -2088
rect 10462 -2140 10514 -2088
rect 11672 -2140 11724 -2088
rect 11882 -2140 11934 -2088
rect 13428 -2726 13480 -2674
rect 1250 -3638 1302 -3586
rect 13428 -3022 13480 -2970
rect 1250 -3880 1302 -3828
rect 1976 -4596 2028 -4544
rect 1785 -4842 1839 -4788
rect 2220 -4596 2272 -4544
rect 2548 -4596 2600 -4544
rect 2774 -4596 2826 -4544
rect 4062 -4596 4114 -4544
rect 4294 -4596 4346 -4544
rect 5584 -4596 5636 -4544
rect 5854 -4596 5906 -4544
rect 7160 -4596 7212 -4544
rect 7450 -4596 7502 -4544
rect 8734 -4596 8786 -4544
rect 8982 -4596 9034 -4544
rect 10322 -4596 10374 -4544
rect 10556 -4596 10608 -4544
rect 11772 -4596 11824 -4544
rect 12010 -4596 12062 -4544
rect 12896 -4596 12948 -4544
rect 2317 -4842 2371 -4788
rect 13468 -3436 13520 -3384
rect 13468 -3676 13520 -3624
rect 13314 -4596 13366 -4544
<< metal2 >>
rect 2246 -2088 2298 -2082
rect 3958 -2088 4010 -2082
rect 5522 -2088 5574 -2082
rect 8640 -2088 8692 -2082
rect 10226 -2088 10278 -2082
rect 11672 -2088 11724 -2082
rect 2720 -2091 2726 -2088
rect 2298 -2137 2726 -2091
rect 2720 -2140 2726 -2137
rect 2778 -2140 2784 -2088
rect 4258 -2091 4264 -2088
rect 4010 -2137 4264 -2091
rect 4258 -2140 4264 -2137
rect 4316 -2140 4322 -2088
rect 5746 -2091 5752 -2088
rect 5574 -2137 5752 -2091
rect 5746 -2140 5752 -2137
rect 5804 -2140 5810 -2088
rect 7106 -2140 7112 -2088
rect 7164 -2091 7170 -2088
rect 7330 -2091 7336 -2088
rect 7164 -2137 7336 -2091
rect 7164 -2140 7170 -2137
rect 7330 -2140 7336 -2137
rect 7388 -2140 7394 -2088
rect 8904 -2091 8910 -2088
rect 8692 -2137 8910 -2091
rect 8904 -2140 8910 -2137
rect 8962 -2140 8968 -2088
rect 10456 -2091 10462 -2088
rect 10278 -2137 10462 -2091
rect 10456 -2140 10462 -2137
rect 10514 -2140 10520 -2088
rect 11876 -2091 11882 -2088
rect 11724 -2137 11882 -2091
rect 11876 -2140 11882 -2137
rect 11934 -2140 11940 -2088
rect 2246 -2146 2298 -2140
rect 3958 -2146 4010 -2140
rect 5522 -2146 5574 -2140
rect 8640 -2146 8692 -2140
rect 10226 -2146 10278 -2140
rect 11672 -2146 11724 -2140
rect 13428 -2674 13480 -2668
rect 13428 -2732 13480 -2726
rect 13436 -2970 13472 -2732
rect 13422 -3022 13428 -2970
rect 13480 -3022 13486 -2970
rect 13468 -3384 13520 -3378
rect 13468 -3442 13520 -3436
rect 1250 -3586 1302 -3580
rect 13475 -3624 13513 -3442
rect 1250 -3644 1302 -3638
rect 1255 -3822 1297 -3644
rect 13462 -3676 13468 -3624
rect 13520 -3676 13526 -3624
rect 1250 -3828 1302 -3822
rect 1250 -3886 1302 -3880
rect 1976 -4544 2028 -4538
rect 2548 -4544 2600 -4538
rect 4062 -4544 4114 -4538
rect 5584 -4544 5636 -4538
rect 7160 -4544 7212 -4538
rect 8734 -4544 8786 -4538
rect 10322 -4544 10374 -4538
rect 11772 -4544 11824 -4538
rect 12896 -4544 12948 -4538
rect 2214 -4546 2220 -4544
rect 2028 -4594 2220 -4546
rect 2214 -4596 2220 -4594
rect 2272 -4596 2278 -4544
rect 2768 -4546 2774 -4544
rect 2600 -4594 2774 -4546
rect 2768 -4596 2774 -4594
rect 2826 -4596 2832 -4544
rect 4288 -4546 4294 -4544
rect 4114 -4594 4294 -4546
rect 4288 -4596 4294 -4594
rect 4346 -4596 4352 -4544
rect 5848 -4546 5854 -4544
rect 5636 -4594 5854 -4546
rect 5848 -4596 5854 -4594
rect 5906 -4596 5912 -4544
rect 7444 -4546 7450 -4544
rect 7212 -4594 7450 -4546
rect 7444 -4596 7450 -4594
rect 7502 -4596 7508 -4544
rect 8976 -4546 8982 -4544
rect 8786 -4594 8982 -4546
rect 8976 -4596 8982 -4594
rect 9034 -4596 9040 -4544
rect 10550 -4546 10556 -4544
rect 10374 -4594 10556 -4546
rect 10550 -4596 10556 -4594
rect 10608 -4596 10614 -4544
rect 12004 -4546 12010 -4544
rect 11824 -4594 12010 -4546
rect 12004 -4596 12010 -4594
rect 12062 -4596 12068 -4544
rect 13308 -4546 13314 -4544
rect 12948 -4594 13314 -4546
rect 13308 -4596 13314 -4594
rect 13366 -4596 13372 -4544
rect 1976 -4602 2028 -4596
rect 2548 -4602 2600 -4596
rect 4062 -4602 4114 -4596
rect 5584 -4602 5636 -4596
rect 7160 -4602 7212 -4596
rect 8734 -4602 8786 -4596
rect 10322 -4602 10374 -4596
rect 11772 -4602 11824 -4596
rect 12896 -4602 12948 -4596
rect 2317 -4788 2371 -4782
rect 1779 -4842 1785 -4788
rect 1839 -4842 2317 -4788
rect 2317 -4848 2371 -4842
use sky130_fd_pr__pfet_01v8_HBKBCU  sky130_fd_pr__pfet_01v8_HBKBCU_0
timestamp 1713286823
transform 1 0 1444 0 1 -3033
box -214 -399 214 399
use cs_inv  x1
timestamp 1713639308
transform 1 0 2117 0 1 -2610
box 293 -2038 1671 576
use cs_inv  x2
timestamp 1713639308
transform 1 0 5157 0 1 -2596
box 293 -2038 1671 576
use cs_inv  x3
timestamp 1713639308
transform 1 0 9837 0 1 -2604
box 293 -2038 1671 576
use cs_inv  x4
timestamp 1713639308
transform 1 0 8319 0 1 -2600
box 293 -2038 1671 576
use cs_inv  x5
timestamp 1713639308
transform 1 0 6757 0 1 -2604
box 293 -2038 1671 576
use cs_inv  x6
timestamp 1713639308
transform 1 0 11315 0 1 -2610
box 293 -2038 1671 576
use cs_inv  x7
timestamp 1713639308
transform 1 0 3635 0 1 -2600
box 293 -2038 1671 576
use sky130_fd_pr__nfet_01v8_6FB46G  XM21
timestamp 1713284121
transform 1 0 1442 0 1 -3858
box -214 -252 214 252
use sky130_fd_pr__nfet_01v8_4BNSKG  XM23
timestamp 1713275267
transform 1 0 13688 0 1 -3640
box -214 -252 214 252
use sky130_fd_pr__pfet_01v8_X4438S  XM24
timestamp 1713275267
transform 1 0 13698 0 1 -3001
box -214 -291 214 291
<< labels >>
flabel metal1 13598 -2680 13798 -2480 0 FreeSans 256 0 0 0 VDD
port 11 nsew
flabel metal1 13592 -4136 13792 -3936 0 FreeSans 256 0 0 0 GND
port 12 nsew
flabel metal1 14054 -3340 14254 -3140 0 FreeSans 256 0 0 0 osc
port 4 nsew
flabel metal1 442 -3980 642 -3780 0 FreeSans 256 0 0 0 vctrl
port 19 nsew
flabel metal1 2052 -3206 2052 -3206 0 FreeSans 320 0 0 0 Vp
flabel metal1 1336 -4350 1536 -4150 0 FreeSans 256 0 0 0 GND
port 3 nsew
flabel metal1 1766 -2418 1966 -2218 0 FreeSans 256 0 0 0 VDD
port 9 nsew
<< end >>
