magic
tech sky130A
magscale 1 2
timestamp 1713286823
<< error_p >>
rect -29 261 29 267
rect -29 227 -17 261
rect -29 221 29 227
rect -29 -227 29 -221
rect -29 -261 -17 -227
rect -29 -267 29 -261
<< nwell >>
rect -214 -399 214 399
<< pmos >>
rect -18 -180 18 180
<< pdiff >>
rect -76 168 -18 180
rect -76 -168 -64 168
rect -30 -168 -18 168
rect -76 -180 -18 -168
rect 18 168 76 180
rect 18 -168 30 168
rect 64 -168 76 168
rect 18 -180 76 -168
<< pdiffc >>
rect -64 -168 -30 168
rect 30 -168 64 168
<< nsubdiff >>
rect -178 329 -82 363
rect 82 329 178 363
rect -178 267 -144 329
rect 144 267 178 329
rect -178 -329 -144 -267
rect 144 -329 178 -267
rect -178 -363 -82 -329
rect 82 -363 178 -329
<< nsubdiffcont >>
rect -82 329 82 363
rect -178 -267 -144 267
rect 144 -267 178 267
rect -82 -363 82 -329
<< poly >>
rect -33 261 33 277
rect -33 227 -17 261
rect 17 227 33 261
rect -33 211 33 227
rect -18 180 18 211
rect -18 -211 18 -180
rect -33 -227 33 -211
rect -33 -261 -17 -227
rect 17 -261 33 -227
rect -33 -277 33 -261
<< polycont >>
rect -17 227 17 261
rect -17 -261 17 -227
<< locali >>
rect -178 267 -144 363
rect 144 267 178 363
rect -33 227 -17 261
rect 17 227 33 261
rect -64 168 -30 184
rect -64 -184 -30 -168
rect 30 168 64 184
rect 30 -184 64 -168
rect -33 -261 -17 -227
rect 17 -261 33 -227
rect -178 -329 -144 -267
rect 144 -329 178 -267
rect -178 -363 -82 -329
rect 82 -363 178 -329
<< viali >>
rect -144 329 -82 363
rect -82 329 82 363
rect 82 329 144 363
rect -17 227 17 261
rect -64 17 -30 151
rect 30 -151 64 -17
rect -17 -261 17 -227
<< metal1 >>
rect -156 363 156 369
rect -156 329 -144 363
rect 144 329 156 363
rect -156 323 156 329
rect -29 261 29 267
rect -29 227 -17 261
rect 17 227 29 261
rect -29 221 29 227
rect -70 151 -24 163
rect -70 17 -64 151
rect -30 17 -24 151
rect -70 5 -24 17
rect 24 -17 70 -5
rect 24 -151 30 -17
rect 64 -151 70 -17
rect 24 -163 70 -151
rect -29 -227 29 -221
rect -29 -261 -17 -227
rect 17 -261 29 -227
rect -29 -267 29 -261
<< properties >>
string FIXED_BBOX -161 -346 161 346
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.8 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
