magic
tech sky130A
magscale 1 2
timestamp 1714564928
<< error_p >>
rect -29 114 29 120
rect -29 80 -17 114
rect -29 74 29 80
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect -29 -120 29 -114
<< pwell >>
rect -214 -252 214 252
<< nmos >>
rect -18 -42 18 42
<< ndiff >>
rect -76 30 -18 42
rect -76 -30 -64 30
rect -30 -30 -18 30
rect -76 -42 -18 -30
rect 18 30 76 42
rect 18 -30 30 30
rect 64 -30 76 30
rect 18 -42 76 -30
<< ndiffc >>
rect -64 -30 -30 30
rect 30 -30 64 30
<< psubdiff >>
rect -178 182 -82 216
rect 82 182 178 216
rect -178 120 -144 182
rect 144 120 178 182
rect -178 -182 -144 -120
rect 144 -182 178 -120
rect -178 -216 -82 -182
rect 82 -216 178 -182
<< psubdiffcont >>
rect -82 182 82 216
rect -178 -120 -144 120
rect 144 -120 178 120
rect -82 -216 82 -182
<< poly >>
rect -33 114 33 130
rect -33 80 -17 114
rect 17 80 33 114
rect -33 64 33 80
rect -18 42 18 64
rect -18 -64 18 -42
rect -33 -80 33 -64
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -33 -130 33 -114
<< polycont >>
rect -17 80 17 114
rect -17 -114 17 -80
<< locali >>
rect -178 182 -82 216
rect 82 182 178 216
rect -178 120 -144 182
rect -33 80 -17 114
rect 17 80 33 114
rect -64 30 -30 46
rect -64 -46 -30 -30
rect 30 30 64 46
rect 30 -46 64 -30
rect -33 -114 -17 -80
rect 17 -114 33 -80
rect -178 -182 -144 -120
rect -178 -216 -82 -182
rect 82 -216 178 -182
<< viali >>
rect 144 120 178 182
rect -17 80 17 114
rect -64 -30 -30 30
rect 30 -30 64 30
rect -17 -114 17 -80
rect 144 -120 178 120
rect 144 -182 178 -120
<< metal1 >>
rect 138 182 184 194
rect -29 114 29 120
rect -29 80 -17 114
rect 17 80 29 114
rect -29 74 29 80
rect -70 30 -24 42
rect -70 -30 -64 30
rect -30 -30 -24 30
rect -70 -42 -24 -30
rect 24 30 70 42
rect 24 -30 30 30
rect 64 -30 70 30
rect 24 -42 70 -30
rect -29 -80 29 -74
rect -29 -114 -17 -80
rect 17 -114 29 -80
rect -29 -120 29 -114
rect 138 -182 144 182
rect 178 -182 184 182
rect 138 -194 184 -182
<< properties >>
string FIXED_BBOX -161 -199 161 199
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 100 viagl 0 viagt 0
<< end >>
