magic
tech sky130A
magscale 1 2
timestamp 1714294046
<< error_p >>
rect -29 1572 29 1578
rect -29 1538 -17 1572
rect -29 1532 29 1538
rect -29 -1538 29 -1532
rect -29 -1572 -17 -1538
rect -29 -1578 29 -1572
<< pwell >>
rect -214 -1710 214 1710
<< nmos >>
rect -18 -1500 18 1500
<< ndiff >>
rect -76 1488 -18 1500
rect -76 -1488 -64 1488
rect -30 -1488 -18 1488
rect -76 -1500 -18 -1488
rect 18 1488 76 1500
rect 18 -1488 30 1488
rect 64 -1488 76 1488
rect 18 -1500 76 -1488
<< ndiffc >>
rect -64 -1488 -30 1488
rect 30 -1488 64 1488
<< psubdiff >>
rect -178 1640 -82 1674
rect 82 1640 178 1674
rect -178 1578 -144 1640
rect 144 1578 178 1640
rect -178 -1640 -144 -1578
rect 144 -1640 178 -1578
rect -178 -1674 -82 -1640
rect 82 -1674 178 -1640
<< psubdiffcont >>
rect -82 1640 82 1674
rect -178 -1578 -144 1578
rect 144 -1578 178 1578
rect -82 -1674 82 -1640
<< poly >>
rect -33 1572 33 1588
rect -33 1538 -17 1572
rect 17 1538 33 1572
rect -33 1522 33 1538
rect -18 1500 18 1522
rect -18 -1522 18 -1500
rect -33 -1538 33 -1522
rect -33 -1572 -17 -1538
rect 17 -1572 33 -1538
rect -33 -1588 33 -1572
<< polycont >>
rect -17 1538 17 1572
rect -17 -1572 17 -1538
<< locali >>
rect -178 1640 -82 1674
rect 82 1640 178 1674
rect -178 1578 -144 1640
rect 144 1578 178 1640
rect -33 1538 -17 1572
rect 17 1538 33 1572
rect -64 1488 -30 1504
rect -64 -1504 -30 -1488
rect 30 1488 64 1504
rect 30 -1504 64 -1488
rect -33 -1572 -17 -1538
rect 17 -1572 33 -1538
rect -178 -1674 -144 -1578
rect 144 -1674 178 -1578
<< viali >>
rect -17 1538 17 1572
rect -64 281 -30 1471
rect 30 -1471 64 -281
rect -17 -1572 17 -1538
rect -144 -1674 -82 -1640
rect -82 -1674 82 -1640
rect 82 -1674 144 -1640
<< metal1 >>
rect -29 1572 29 1578
rect -29 1538 -17 1572
rect 17 1538 29 1572
rect -29 1532 29 1538
rect -70 1471 -24 1483
rect -70 281 -64 1471
rect -30 281 -24 1471
rect -70 269 -24 281
rect 24 -281 70 -269
rect 24 -1471 30 -281
rect 64 -1471 70 -281
rect 24 -1483 70 -1471
rect -29 -1538 29 -1532
rect -29 -1572 -17 -1538
rect 17 -1572 29 -1538
rect -29 -1578 29 -1572
rect -156 -1640 156 -1634
rect -156 -1674 -144 -1640
rect 144 -1674 156 -1640
rect -156 -1680 156 -1674
<< properties >>
string FIXED_BBOX -161 -1657 161 1657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 15.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 100 viagr 0 viagl 0 viagt 0
<< end >>
