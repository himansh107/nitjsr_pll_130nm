magic
tech sky130A
magscale 1 2
timestamp 1713639308
<< viali >>
rect 977 266 1175 318
rect 991 -1818 1181 -1784
<< metal1 >>
rect 975 430 1175 576
rect 799 316 805 368
rect 857 366 863 368
rect 913 366 1259 430
rect 857 318 1259 366
rect 857 316 863 318
rect 913 266 977 318
rect 1175 266 1259 318
rect 913 254 1259 266
rect 753 154 1105 184
rect 421 68 621 140
rect 755 68 793 154
rect 1189 96 1195 105
rect 421 14 793 68
rect 421 -60 621 14
rect 755 -86 793 14
rect 859 66 911 72
rect 911 16 1047 64
rect 1109 62 1195 96
rect 1189 53 1195 62
rect 1247 53 1253 105
rect 859 8 911 14
rect 755 -116 1113 -86
rect 613 -420 1109 -372
rect 619 -508 663 -420
rect 533 -564 665 -508
rect 917 -552 923 -500
rect 975 -512 981 -500
rect 975 -540 1041 -512
rect 975 -552 981 -540
rect 1303 -558 1339 -557
rect 293 -784 493 -724
rect 533 -784 589 -564
rect 619 -644 663 -564
rect 1107 -592 1341 -558
rect 619 -692 1115 -644
rect 1303 -750 1339 -592
rect 1471 -750 1671 -670
rect 293 -840 589 -784
rect 1301 -794 1671 -750
rect 293 -924 493 -840
rect 531 -1070 587 -840
rect 859 -938 865 -886
rect 917 -894 923 -886
rect 1303 -894 1339 -794
rect 1471 -870 1671 -794
rect 917 -930 1339 -894
rect 917 -938 923 -930
rect 1303 -934 1339 -930
rect 619 -1044 1115 -996
rect 619 -1070 657 -1044
rect 531 -1126 657 -1070
rect 619 -1192 657 -1126
rect 865 -1084 917 -1078
rect 917 -1094 1019 -1092
rect 917 -1128 1049 -1094
rect 981 -1130 1049 -1128
rect 865 -1142 917 -1136
rect 1111 -1150 1341 -1116
rect 619 -1240 1115 -1192
rect 879 -1464 885 -1412
rect 937 -1421 943 -1412
rect 1306 -1421 1340 -1150
rect 937 -1455 1340 -1421
rect 937 -1464 943 -1455
rect 483 -1550 683 -1504
rect 743 -1536 1115 -1492
rect 743 -1550 787 -1536
rect 483 -1594 787 -1550
rect 483 -1704 683 -1594
rect 741 -1680 785 -1594
rect 879 -1632 885 -1580
rect 937 -1589 943 -1580
rect 937 -1595 1032 -1589
rect 937 -1623 1048 -1595
rect 937 -1632 943 -1623
rect 995 -1629 1048 -1623
rect 1115 -1634 1253 -1600
rect 741 -1724 1111 -1680
rect 1214 -1764 1248 -1634
rect 923 -1784 1249 -1764
rect 923 -1818 991 -1784
rect 1181 -1818 1249 -1784
rect 923 -1852 1249 -1818
rect 985 -2014 1185 -1852
<< via1 >>
rect 805 316 857 368
rect 859 14 911 66
rect 1195 53 1247 105
rect 923 -552 975 -500
rect 865 -938 917 -886
rect 865 -1136 917 -1084
rect 885 -1464 937 -1412
rect 885 -1632 937 -1580
<< metal2 >>
rect 805 368 857 374
rect 805 310 857 316
rect 807 66 855 310
rect 1195 105 1247 111
rect 807 16 859 66
rect 853 14 859 16
rect 911 14 917 66
rect 1195 47 1247 53
rect 1204 -196 1238 47
rect 935 -224 1238 -196
rect 935 -494 963 -224
rect 1204 -227 1238 -224
rect 923 -500 975 -494
rect 923 -558 975 -552
rect 865 -886 917 -880
rect 865 -944 917 -938
rect 873 -1084 909 -944
rect 859 -1136 865 -1084
rect 917 -1136 923 -1084
rect 885 -1412 937 -1406
rect 885 -1470 937 -1464
rect 894 -1574 928 -1470
rect 885 -1580 937 -1574
rect 885 -1638 937 -1632
use sky130_fd_pr__nfet_01v8_4BNSKG  XM1
timestamp 1713275267
transform 1 0 1081 0 1 -1120
box -214 -252 214 252
use sky130_fd_pr__pfet_01v8_X4438S  XM2
timestamp 1713275267
transform 1 0 1079 0 1 35
box -214 -291 214 291
use sky130_fd_pr__pfet_01v8_X4438S  XM3
timestamp 1713275267
transform 1 0 1079 0 1 -529
box -214 -291 214 291
use sky130_fd_pr__nfet_01v8_4BNSKG  XM4
timestamp 1713275267
transform 1 0 1083 0 1 -1606
box -214 -252 214 252
<< labels >>
flabel metal1 421 -60 621 140 0 FreeSans 256 0 0 0 Vp
port 1 nsew
flabel metal1 483 -1704 683 -1504 0 FreeSans 256 0 0 0 Vn
port 4 nsew
flabel metal1 293 -924 493 -724 0 FreeSans 256 0 0 0 in
port 3 nsew
flabel metal1 1471 -870 1671 -670 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 975 376 1175 576 0 FreeSans 256 0 0 0 VDD
port 5 nsew
flabel space 985 -2038 1185 -1838 0 FreeSans 256 0 0 0 GND
port 5 nsew
<< end >>
