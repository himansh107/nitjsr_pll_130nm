magic
tech sky130A
magscale 1 2
timestamp 1714285468
<< error_p >>
rect -29 135 29 141
rect -29 101 -17 135
rect -29 95 29 101
rect -29 -101 29 -95
rect -29 -135 -17 -101
rect -29 -141 29 -135
<< nwell >>
rect -214 -273 214 273
<< pmos >>
rect -18 -54 18 54
<< pdiff >>
rect -76 42 -18 54
rect -76 -42 -64 42
rect -30 -42 -18 42
rect -76 -54 -18 -42
rect 18 42 76 54
rect 18 -42 30 42
rect 64 -42 76 42
rect 18 -54 76 -42
<< pdiffc >>
rect -64 -42 -30 42
rect 30 -42 64 42
<< nsubdiff >>
rect -178 203 -82 237
rect 82 203 178 237
rect -178 141 -144 203
rect 144 141 178 203
rect -178 -203 -144 -141
rect 144 -203 178 -141
rect -178 -237 -82 -203
rect 82 -237 178 -203
<< nsubdiffcont >>
rect -82 203 82 237
rect -178 -141 -144 141
rect 144 -141 178 141
rect -82 -237 82 -203
<< poly >>
rect -33 135 33 151
rect -33 101 -17 135
rect 17 101 33 135
rect -33 85 33 101
rect -18 54 18 85
rect -18 -85 18 -54
rect -33 -101 33 -85
rect -33 -135 -17 -101
rect 17 -135 33 -101
rect -33 -151 33 -135
<< polycont >>
rect -17 101 17 135
rect -17 -135 17 -101
<< locali >>
rect -178 203 -82 237
rect 82 203 178 237
rect -178 141 -144 203
rect -33 101 -17 135
rect 17 101 33 135
rect -64 42 -30 58
rect -64 -58 -30 -42
rect 30 42 64 58
rect 30 -58 64 -42
rect -33 -135 -17 -101
rect 17 -135 33 -101
rect -178 -203 -144 -141
rect -178 -237 -82 -203
rect 82 -237 178 -203
<< viali >>
rect 144 141 178 203
rect -17 101 17 135
rect -64 -42 -30 42
rect 30 -42 64 42
rect -17 -135 17 -101
rect 144 -141 178 141
rect 144 -203 178 -141
<< metal1 >>
rect 138 203 184 215
rect -29 135 29 141
rect -29 101 -17 135
rect 17 101 29 135
rect -29 95 29 101
rect -70 42 -24 54
rect -70 -42 -64 42
rect -30 -42 -24 42
rect -70 -54 -24 -42
rect 24 42 70 54
rect 24 -42 30 42
rect 64 -42 70 42
rect 24 -54 70 -42
rect -29 -101 29 -95
rect -29 -135 -17 -101
rect 17 -135 29 -101
rect -29 -141 29 -135
rect 138 -203 144 203
rect 178 -203 184 203
rect 138 -215 184 -203
<< properties >>
string FIXED_BBOX -161 -220 161 220
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.54 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 100 viagl 0 viagt 0
<< end >>
