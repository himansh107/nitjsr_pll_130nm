VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.975 0.995 2.215 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.145 0.995 1.455 1.325 ;
        RECT 1.145 0.825 1.350 0.995 ;
        RECT 1.000 0.300 1.350 0.825 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.995 0.975 1.325 ;
        RECT 0.595 0.300 0.810 0.995 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.995 0.395 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.085 0.425 0.825 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.295 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.915 1.835 2.195 2.635 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.385 1.665 1.715 2.465 ;
        RECT 0.515 1.495 1.795 1.665 ;
        RECT 1.625 0.825 1.795 1.495 ;
        RECT 1.520 0.255 2.215 0.825 ;
    END
  END Y
END sky130_fd_sc_hd__nand4_1
MACRO sky130_fd_sc_hd__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.755 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.765 1.240 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.745 0.330 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.085 0.345 0.575 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.245 2.635 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.415 1.665 1.745 2.465 ;
        RECT 0.515 1.495 1.745 1.665 ;
        RECT 0.515 0.595 0.695 1.495 ;
        RECT 1.415 0.595 1.745 0.825 ;
        RECT 0.515 0.255 1.745 0.595 ;
    END
  END Y
END sky130_fd_sc_hd__nand3_1
MACRO sky130_fd_sc_hd__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvpwrvgnd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER li1 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.085 1.470 0.375 2.635 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
END sky130_fd_sc_hd__tapvpwrvgnd_1
MACRO sky130_fd_sc_hd__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.320 1.075 0.650 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.320 0.085 0.550 0.905 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.210 0.105 1.140 1.015 ;
        RECT 0.210 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.340 1.495 0.550 2.635 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.720 1.485 1.050 2.465 ;
        RECT 0.820 0.885 1.050 1.485 ;
        RECT 0.720 0.255 1.050 0.885 ;
    END
  END Y
END sky130_fd_sc_hd__inv_1
MACRO sky130_fd_sc_hd__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.940 1.075 1.275 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.430 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.085 0.395 0.885 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.105 1.375 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.085 1.495 0.365 2.635 ;
        RECT 1.035 1.495 1.295 2.635 ;
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.485 0.865 2.465 ;
        RECT 0.600 0.885 0.770 1.485 ;
        RECT 0.600 0.255 1.295 0.885 ;
    END
  END Y
END sky130_fd_sc_hd__nand2_1
MACRO pfd_lay
  CLASS BLOCK ;
  FOREIGN pfd_lay ;
  ORIGIN -3.250 15.880 ;
  SIZE 28.700 BY 22.490 ;
  PIN f_clk_in
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 6.950 2.900 7.280 2.915 ;
        RECT 5.950 2.700 7.280 2.900 ;
        RECT 6.950 2.675 7.280 2.700 ;
      LAYER met1 ;
        RECT 4.250 2.900 5.250 3.380 ;
        RECT 5.920 2.900 6.180 2.960 ;
        RECT 4.250 2.700 6.180 2.900 ;
        RECT 4.250 2.380 5.250 2.700 ;
        RECT 5.920 2.640 6.180 2.700 ;
    END
  END f_clk_in
  PIN up
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 26.210 3.085 26.540 4.065 ;
        RECT 26.310 2.900 26.540 3.085 ;
        RECT 26.310 2.700 27.950 2.900 ;
        RECT 26.310 2.485 26.540 2.700 ;
        RECT 26.210 1.855 26.540 2.485 ;
      LAYER met1 ;
        RECT 27.670 2.900 27.930 2.960 ;
        RECT 28.800 2.900 29.800 3.300 ;
        RECT 27.670 2.700 29.800 2.900 ;
        RECT 27.670 2.640 27.930 2.700 ;
        RECT 28.800 2.300 29.800 2.700 ;
    END
  END up
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 13.120 -0.655 14.880 -0.605 ;
        RECT 9.270 -0.660 11.300 -0.655 ;
        RECT 12.570 -0.660 14.880 -0.655 ;
        RECT 9.270 -0.675 14.880 -0.660 ;
        RECT 8.630 -2.210 14.880 -0.675 ;
        RECT 8.630 -2.260 13.580 -2.210 ;
        RECT 8.630 -2.280 9.470 -2.260 ;
      LAYER li1 ;
        RECT 8.905 -2.005 9.195 -0.840 ;
        RECT 9.545 -1.985 9.825 -0.845 ;
        RECT 10.495 -1.985 10.755 -0.845 ;
        RECT 13.395 -1.935 13.675 -0.795 ;
        RECT 14.345 -1.935 14.605 -0.795 ;
        RECT 8.820 -2.175 9.280 -2.005 ;
        RECT 9.460 -2.155 10.840 -1.985 ;
        RECT 13.310 -2.105 14.690 -1.935 ;
      LAYER met1 ;
        RECT 8.820 -2.040 9.280 -1.850 ;
        RECT 9.460 -2.040 10.840 -1.830 ;
        RECT 13.310 -2.040 14.690 -1.780 ;
        RECT 8.820 -2.330 15.180 -2.040 ;
        RECT 9.200 -2.720 15.180 -2.330 ;
        RECT 12.420 -3.400 13.420 -2.720 ;
    END
    PORT
      LAYER nwell ;
        RECT 27.890 -8.410 28.730 -8.400 ;
        RECT 7.360 -10.005 28.730 -8.410 ;
        RECT 7.360 -10.015 27.980 -10.005 ;
      LAYER li1 ;
        RECT 7.550 -8.685 8.930 -8.515 ;
        RECT 11.230 -8.685 12.610 -8.515 ;
        RECT 15.370 -8.685 16.750 -8.515 ;
        RECT 18.590 -8.685 19.970 -8.515 ;
        RECT 22.270 -8.685 24.110 -8.515 ;
        RECT 26.410 -8.685 27.790 -8.515 ;
        RECT 28.080 -8.675 28.540 -8.505 ;
        RECT 7.890 -9.825 8.100 -8.685 ;
        RECT 11.315 -9.825 11.595 -8.685 ;
        RECT 12.265 -9.825 12.525 -8.685 ;
        RECT 15.710 -9.825 15.920 -8.685 ;
        RECT 18.930 -9.825 19.140 -8.685 ;
        RECT 22.360 -9.825 22.615 -8.685 ;
        RECT 23.285 -9.485 23.515 -8.685 ;
        RECT 26.750 -9.825 26.960 -8.685 ;
        RECT 28.165 -9.840 28.455 -8.675 ;
      LAYER met1 ;
        RECT 17.940 -8.025 18.940 -7.160 ;
        RECT 7.830 -8.160 27.970 -8.025 ;
        RECT 7.830 -8.350 28.520 -8.160 ;
        RECT 7.830 -8.360 28.540 -8.350 ;
        RECT 7.550 -8.830 28.540 -8.360 ;
        RECT 7.550 -8.840 28.150 -8.830 ;
        RECT 7.830 -8.845 28.150 -8.840 ;
        RECT 27.900 -8.850 28.150 -8.845 ;
    END
    PORT
      LAYER nwell ;
        RECT 10.580 -13.075 14.550 -13.015 ;
        RECT 10.580 -13.145 15.570 -13.075 ;
        RECT 10.580 -14.620 16.240 -13.145 ;
        RECT 13.810 -14.680 16.240 -14.620 ;
        RECT 15.400 -14.750 16.240 -14.680 ;
      LAYER li1 ;
        RECT 10.855 -14.345 11.115 -13.205 ;
        RECT 11.785 -14.345 12.065 -13.205 ;
        RECT 10.770 -14.515 12.150 -14.345 ;
        RECT 14.085 -14.405 14.345 -13.265 ;
        RECT 15.015 -14.405 15.295 -13.265 ;
        RECT 14.000 -14.575 15.380 -14.405 ;
        RECT 15.675 -14.475 15.965 -13.310 ;
        RECT 15.590 -14.645 16.050 -14.475 ;
      LAYER met1 ;
        RECT 10.770 -14.620 12.150 -14.190 ;
        RECT 14.000 -14.620 15.380 -14.250 ;
        RECT 15.590 -14.620 16.050 -14.320 ;
        RECT 10.580 -14.800 16.050 -14.620 ;
        RECT 10.580 -14.960 15.640 -14.800 ;
        RECT 13.340 -15.880 14.340 -14.960 ;
    END
    PORT
      LAYER nwell ;
        RECT 19.900 -2.905 23.660 -1.300 ;
      LAYER li1 ;
        RECT 20.090 -1.575 22.390 -1.405 ;
        RECT 23.010 -1.575 23.470 -1.405 ;
        RECT 20.175 -2.715 20.435 -1.575 ;
        RECT 21.105 -2.375 21.275 -1.575 ;
        RECT 22.005 -2.375 22.285 -1.575 ;
        RECT 23.095 -2.740 23.385 -1.575 ;
      LAYER met1 ;
        RECT 20.800 -1.250 21.800 -0.500 ;
        RECT 20.090 -1.730 23.470 -1.250 ;
        RECT 22.250 -1.750 23.220 -1.730 ;
    END
    PORT
      LAYER nwell ;
        RECT 6.440 2.905 27.520 4.510 ;
      LAYER li1 ;
        RECT 6.630 4.235 8.010 4.405 ;
        RECT 10.310 4.235 11.690 4.405 ;
        RECT 14.450 4.235 15.830 4.405 ;
        RECT 17.670 4.235 19.050 4.405 ;
        RECT 21.350 4.235 23.190 4.405 ;
        RECT 25.490 4.235 27.330 4.405 ;
        RECT 6.970 3.095 7.180 4.235 ;
        RECT 10.395 3.095 10.675 4.235 ;
        RECT 11.345 3.095 11.605 4.235 ;
        RECT 14.790 3.095 15.000 4.235 ;
        RECT 18.010 3.095 18.220 4.235 ;
        RECT 21.440 3.095 21.695 4.235 ;
        RECT 22.365 3.435 22.595 4.235 ;
        RECT 25.830 3.095 26.040 4.235 ;
        RECT 26.955 3.070 27.245 4.235 ;
      LAYER met1 ;
        RECT 16.560 5.240 17.560 6.100 ;
        RECT 6.900 4.760 27.040 5.240 ;
        RECT 6.900 4.560 27.600 4.760 ;
        RECT 6.630 4.420 27.600 4.560 ;
        RECT 6.630 4.080 8.010 4.420 ;
        RECT 10.310 4.080 11.690 4.420 ;
        RECT 14.450 4.080 15.830 4.420 ;
        RECT 17.670 4.080 19.050 4.420 ;
        RECT 21.350 4.080 23.190 4.420 ;
        RECT 25.490 4.080 27.330 4.420 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 28.095 -11.120 28.525 -10.335 ;
        RECT 15.605 -12.815 16.035 -12.030 ;
      LAYER li1 ;
        RECT 7.870 -11.235 8.100 -10.415 ;
        RECT 11.315 -11.235 11.625 -10.435 ;
        RECT 15.690 -11.235 15.920 -10.415 ;
        RECT 18.910 -11.235 19.140 -10.415 ;
        RECT 22.360 -11.235 22.615 -10.745 ;
        RECT 26.730 -11.235 26.960 -10.415 ;
        RECT 28.165 -11.225 28.455 -10.500 ;
        RECT 7.550 -11.405 8.930 -11.235 ;
        RECT 11.230 -11.405 12.610 -11.235 ;
        RECT 15.370 -11.405 16.750 -11.235 ;
        RECT 18.590 -11.405 19.970 -11.235 ;
        RECT 22.270 -11.405 24.110 -11.235 ;
        RECT 26.410 -11.405 27.790 -11.235 ;
        RECT 28.080 -11.395 28.540 -11.225 ;
        RECT 10.770 -11.795 12.150 -11.625 ;
        RECT 11.755 -12.595 12.065 -11.795 ;
        RECT 14.000 -11.855 15.380 -11.685 ;
        RECT 14.985 -12.655 15.295 -11.855 ;
        RECT 15.590 -11.925 16.050 -11.755 ;
        RECT 15.675 -12.650 15.965 -11.925 ;
      LAYER met1 ;
        RECT 27.900 -11.070 28.200 -11.050 ;
        RECT 27.900 -11.080 28.540 -11.070 ;
        RECT 7.550 -11.220 28.540 -11.080 ;
        RECT 7.360 -11.550 28.540 -11.220 ;
        RECT 7.360 -11.560 28.520 -11.550 ;
        RECT 7.360 -11.900 28.010 -11.560 ;
        RECT 10.770 -11.950 12.150 -11.900 ;
        RECT 14.000 -12.010 15.380 -11.900 ;
        RECT 15.590 -12.080 16.050 -11.900 ;
        RECT 25.000 -12.400 26.000 -11.900 ;
    END
    PORT
      LAYER pwell ;
        RECT 23.025 -4.020 23.455 -3.235 ;
      LAYER li1 ;
        RECT 20.180 -4.125 20.515 -3.385 ;
        RECT 23.095 -4.125 23.385 -3.400 ;
        RECT 20.090 -4.295 22.390 -4.125 ;
        RECT 23.010 -4.295 23.470 -4.125 ;
      LAYER met1 ;
        RECT 22.250 -3.970 23.220 -3.950 ;
        RECT 20.090 -4.450 23.470 -3.970 ;
        RECT 21.350 -5.250 22.350 -4.450 ;
    END
    PORT
      LAYER pwell ;
        RECT 26.885 1.790 27.315 2.575 ;
        RECT 8.835 -0.345 9.265 0.440 ;
      LAYER li1 ;
        RECT 6.950 1.685 7.180 2.505 ;
        RECT 10.395 1.685 10.705 2.485 ;
        RECT 14.770 1.685 15.000 2.505 ;
        RECT 17.990 1.685 18.220 2.505 ;
        RECT 21.440 1.685 21.695 2.175 ;
        RECT 25.810 1.685 26.040 2.505 ;
        RECT 26.955 1.685 27.245 2.410 ;
        RECT 6.630 1.515 8.010 1.685 ;
        RECT 10.310 1.515 11.690 1.685 ;
        RECT 14.450 1.515 15.830 1.685 ;
        RECT 17.670 1.515 19.050 1.685 ;
        RECT 21.350 1.515 23.190 1.685 ;
        RECT 25.490 1.515 27.330 1.685 ;
        RECT 8.820 0.545 9.280 0.715 ;
        RECT 9.460 0.565 10.840 0.735 ;
        RECT 13.310 0.615 14.690 0.785 ;
        RECT 8.905 -0.180 9.195 0.545 ;
        RECT 9.545 -0.235 9.855 0.565 ;
        RECT 13.395 -0.185 13.705 0.615 ;
      LAYER met1 ;
        RECT 6.630 1.500 8.010 1.840 ;
        RECT 10.310 1.500 11.690 1.840 ;
        RECT 14.450 1.500 15.830 1.840 ;
        RECT 17.670 1.500 19.050 1.840 ;
        RECT 21.350 1.500 23.190 1.840 ;
        RECT 25.490 1.500 27.330 1.840 ;
        RECT 6.630 1.360 27.330 1.500 ;
        RECT 6.900 1.020 27.600 1.360 ;
        RECT 6.900 0.680 27.040 1.020 ;
        RECT 8.820 0.390 9.280 0.680 ;
        RECT 9.460 0.410 10.840 0.680 ;
        RECT 13.310 0.460 14.690 0.680 ;
        RECT 17.020 0.000 18.020 0.680 ;
    END
  END VGND
  PIN down
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 27.130 -9.835 27.460 -8.855 ;
        RECT 27.230 -10.050 27.460 -9.835 ;
        RECT 27.230 -10.250 29.900 -10.050 ;
        RECT 27.230 -10.435 27.460 -10.250 ;
        RECT 27.130 -11.065 27.460 -10.435 ;
      LAYER met1 ;
        RECT 29.670 -10.050 29.930 -9.990 ;
        RECT 30.950 -10.050 31.950 -9.500 ;
        RECT 29.670 -10.250 31.950 -10.050 ;
        RECT 29.670 -10.310 29.930 -10.250 ;
        RECT 30.950 -10.500 31.950 -10.250 ;
    END
  END down
  PIN f_vco
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 6.900 -10.005 8.170 -10.000 ;
        RECT 6.900 -10.200 8.200 -10.005 ;
        RECT 7.870 -10.245 8.200 -10.200 ;
      LAYER met1 ;
        RECT 3.250 -10.000 4.250 -9.700 ;
        RECT 4.820 -10.000 5.080 -9.940 ;
        RECT 3.250 -10.200 5.080 -10.000 ;
        RECT 3.250 -10.700 4.250 -10.200 ;
        RECT 4.820 -10.260 5.080 -10.200 ;
        RECT 6.190 -10.000 6.510 -9.970 ;
        RECT 6.870 -10.000 7.130 -9.940 ;
        RECT 6.190 -10.200 7.130 -10.000 ;
        RECT 6.190 -10.230 6.510 -10.200 ;
        RECT 6.870 -10.260 7.130 -10.200 ;
      LAYER met2 ;
        RECT 4.790 -10.000 5.110 -9.970 ;
        RECT 6.220 -10.000 6.480 -9.940 ;
        RECT 4.790 -10.200 6.480 -10.000 ;
        RECT 4.790 -10.230 5.110 -10.200 ;
        RECT 6.220 -10.260 6.480 -10.200 ;
    END
  END VPWR
  OBS
      LAYER pwell ;
        RECT 6.840 1.705 7.770 2.615 ;
        RECT 10.335 1.705 11.685 2.615 ;
        RECT 14.660 1.705 15.590 2.615 ;
        RECT 17.880 1.705 18.810 2.615 ;
        RECT 21.355 1.705 23.185 2.615 ;
        RECT 25.700 1.705 26.630 2.615 ;
        RECT 6.840 1.685 6.945 1.705 ;
        RECT 6.775 1.515 6.945 1.685 ;
        RECT 10.450 1.515 10.620 1.705 ;
        RECT 14.660 1.685 14.765 1.705 ;
        RECT 17.880 1.685 17.985 1.705 ;
        RECT 14.595 1.515 14.765 1.685 ;
        RECT 17.815 1.515 17.985 1.685 ;
        RECT 21.500 1.515 21.670 1.705 ;
        RECT 25.700 1.685 25.805 1.705 ;
        RECT 25.635 1.515 25.805 1.685 ;
        RECT 9.600 0.545 9.770 0.735 ;
        RECT 13.450 0.595 13.620 0.785 ;
        RECT 9.485 -0.365 10.835 0.545 ;
        RECT 13.335 -0.315 14.685 0.595 ;
        RECT 20.095 -4.105 22.385 -3.195 ;
        RECT 20.240 -4.295 20.410 -4.105 ;
        RECT 7.760 -11.215 8.690 -10.305 ;
        RECT 11.255 -11.215 12.605 -10.305 ;
        RECT 15.580 -11.215 16.510 -10.305 ;
        RECT 18.800 -11.215 19.730 -10.305 ;
        RECT 22.275 -11.215 24.105 -10.305 ;
        RECT 26.620 -11.215 27.550 -10.305 ;
        RECT 7.760 -11.235 7.865 -11.215 ;
        RECT 7.695 -11.405 7.865 -11.235 ;
        RECT 11.370 -11.405 11.540 -11.215 ;
        RECT 15.580 -11.235 15.685 -11.215 ;
        RECT 18.800 -11.235 18.905 -11.215 ;
        RECT 15.515 -11.405 15.685 -11.235 ;
        RECT 18.735 -11.405 18.905 -11.235 ;
        RECT 22.420 -11.405 22.590 -11.215 ;
        RECT 26.620 -11.235 26.725 -11.215 ;
        RECT 26.555 -11.405 26.725 -11.235 ;
        RECT 11.840 -11.815 12.010 -11.625 ;
        RECT 10.775 -12.725 12.125 -11.815 ;
        RECT 15.070 -11.875 15.240 -11.685 ;
        RECT 14.005 -12.785 15.355 -11.875 ;
      LAYER li1 ;
        RECT 7.350 3.085 7.680 4.065 ;
        RECT 10.845 3.085 11.175 4.065 ;
        RECT 13.175 3.475 13.925 3.730 ;
        RECT 7.450 2.900 7.680 3.085 ;
        RECT 10.405 2.900 10.740 2.925 ;
        RECT 7.450 2.700 10.740 2.900 ;
        RECT 7.450 2.485 7.680 2.700 ;
        RECT 10.405 2.655 10.740 2.700 ;
        RECT 7.350 1.855 7.680 2.485 ;
        RECT 10.910 2.485 11.080 3.085 ;
        RECT 11.250 2.900 11.585 2.925 ;
        RECT 13.700 2.900 13.890 3.475 ;
        RECT 15.170 3.085 15.500 4.065 ;
        RECT 18.390 3.085 18.720 4.065 ;
        RECT 14.770 2.900 15.100 2.915 ;
        RECT 11.250 2.700 12.350 2.900 ;
        RECT 13.700 2.700 15.100 2.900 ;
        RECT 11.250 2.675 11.585 2.700 ;
        RECT 10.910 2.200 11.605 2.485 ;
        RECT 13.700 2.200 13.900 2.700 ;
        RECT 14.770 2.675 15.100 2.700 ;
        RECT 15.270 2.900 15.500 3.085 ;
        RECT 17.990 2.900 18.320 2.915 ;
        RECT 15.270 2.700 18.320 2.900 ;
        RECT 15.270 2.485 15.500 2.700 ;
        RECT 17.990 2.675 18.320 2.700 ;
        RECT 18.490 2.850 18.720 3.085 ;
        RECT 19.900 2.850 20.100 3.800 ;
        RECT 21.865 3.265 22.195 4.065 ;
        RECT 22.765 3.265 23.095 4.065 ;
        RECT 21.865 3.095 23.095 3.265 ;
        RECT 24.400 3.250 25.050 3.450 ;
        RECT 21.460 2.850 21.680 2.925 ;
        RECT 18.490 2.650 20.100 2.850 ;
        RECT 20.750 2.650 21.680 2.850 ;
        RECT 18.490 2.485 18.720 2.650 ;
        RECT 10.910 2.000 13.900 2.200 ;
        RECT 10.910 1.855 11.605 2.000 ;
        RECT 15.170 1.855 15.500 2.485 ;
        RECT 18.390 1.855 18.720 2.485 ;
        RECT 20.750 1.800 20.950 2.650 ;
        RECT 21.460 2.345 21.680 2.650 ;
        RECT 21.865 2.195 22.045 3.095 ;
        RECT 22.215 2.365 22.590 2.925 ;
        RECT 22.795 2.900 23.105 2.925 ;
        RECT 24.850 2.900 25.050 3.250 ;
        RECT 25.810 2.900 26.140 2.915 ;
        RECT 22.795 2.650 24.100 2.900 ;
        RECT 24.850 2.700 26.140 2.900 ;
        RECT 22.795 2.595 23.105 2.650 ;
        RECT 22.765 2.195 23.095 2.425 ;
        RECT 23.855 2.405 24.050 2.650 ;
        RECT 21.865 2.150 23.095 2.195 ;
        RECT 24.850 2.150 25.050 2.700 ;
        RECT 25.810 2.675 26.140 2.700 ;
        RECT 21.865 1.950 25.050 2.150 ;
        RECT 21.865 1.855 23.095 1.950 ;
        RECT 10.060 0.250 10.755 0.395 ;
        RECT 10.060 0.050 11.750 0.250 ;
        RECT 13.910 0.200 14.605 0.445 ;
        RECT 10.060 -0.235 10.755 0.050 ;
        RECT 13.910 0.000 15.900 0.200 ;
        RECT 13.910 -0.185 14.605 0.000 ;
        RECT 9.555 -0.450 9.890 -0.405 ;
        RECT 8.400 -0.650 9.890 -0.450 ;
        RECT 9.555 -0.675 9.890 -0.650 ;
        RECT 10.060 -0.835 10.230 -0.235 ;
        RECT 13.405 -0.400 13.740 -0.355 ;
        RECT 10.400 -0.450 10.735 -0.425 ;
        RECT 10.400 -0.650 12.350 -0.450 ;
        RECT 12.650 -0.600 13.740 -0.400 ;
        RECT 13.405 -0.625 13.740 -0.600 ;
        RECT 10.400 -0.675 10.735 -0.650 ;
        RECT 9.995 -1.815 10.325 -0.835 ;
        RECT 11.425 -0.950 11.625 -0.650 ;
        RECT 13.910 -0.785 14.080 -0.185 ;
        RECT 14.250 -0.415 14.585 -0.375 ;
        RECT 14.250 -0.585 15.185 -0.415 ;
        RECT 14.250 -0.625 14.585 -0.585 ;
        RECT 13.845 -1.765 14.175 -0.785 ;
        RECT 18.600 -2.250 18.800 -1.600 ;
        RECT 18.600 -2.450 19.550 -2.250 ;
        RECT 20.605 -2.545 20.935 -1.745 ;
        RECT 21.475 -2.545 21.805 -1.745 ;
        RECT 20.605 -2.715 21.885 -2.545 ;
        RECT 17.640 -2.950 19.760 -2.940 ;
        RECT 20.200 -2.950 20.485 -2.885 ;
        RECT 17.640 -3.150 20.500 -2.950 ;
        RECT 17.640 -3.160 19.760 -3.150 ;
        RECT 20.200 -3.215 20.485 -3.150 ;
        RECT 20.685 -3.215 21.065 -2.885 ;
        RECT 21.235 -3.215 21.545 -2.885 ;
        RECT 18.700 -3.800 19.800 -3.600 ;
        RECT 18.705 -5.145 18.895 -3.800 ;
        RECT 20.685 -3.910 20.900 -3.215 ;
        RECT 21.235 -3.385 21.440 -3.215 ;
        RECT 21.715 -3.385 21.885 -2.715 ;
        RECT 22.065 -2.950 22.305 -2.545 ;
        RECT 22.065 -3.150 24.850 -2.950 ;
        RECT 22.065 -3.215 22.305 -3.150 ;
        RECT 21.090 -3.910 21.440 -3.385 ;
        RECT 21.610 -3.955 22.305 -3.385 ;
        RECT 8.270 -9.835 8.600 -8.855 ;
        RECT 11.765 -9.835 12.095 -8.855 ;
        RECT 16.090 -9.835 16.420 -8.855 ;
        RECT 19.310 -9.835 19.640 -8.855 ;
        RECT 8.370 -10.050 8.600 -9.835 ;
        RECT 11.325 -10.050 11.660 -9.995 ;
        RECT 8.370 -10.250 11.660 -10.050 ;
        RECT 8.370 -10.435 8.600 -10.250 ;
        RECT 11.325 -10.265 11.660 -10.250 ;
        RECT 8.270 -11.065 8.600 -10.435 ;
        RECT 11.830 -10.435 12.000 -9.835 ;
        RECT 12.170 -10.000 12.505 -9.995 ;
        RECT 16.190 -10.000 16.420 -9.835 ;
        RECT 12.170 -10.200 13.250 -10.000 ;
        RECT 14.850 -10.005 15.950 -10.000 ;
        RECT 16.190 -10.005 19.150 -10.000 ;
        RECT 14.850 -10.200 16.020 -10.005 ;
        RECT 12.170 -10.245 12.505 -10.200 ;
        RECT 11.830 -10.700 12.525 -10.435 ;
        RECT 14.200 -10.700 14.400 -10.250 ;
        RECT 14.850 -10.700 15.050 -10.200 ;
        RECT 15.690 -10.245 16.020 -10.200 ;
        RECT 16.190 -10.200 19.240 -10.005 ;
        RECT 16.190 -10.435 16.420 -10.200 ;
        RECT 18.910 -10.245 19.240 -10.200 ;
        RECT 19.410 -10.050 19.640 -9.835 ;
        RECT 22.785 -9.655 23.115 -8.855 ;
        RECT 23.685 -9.655 24.015 -8.855 ;
        RECT 22.785 -9.825 24.015 -9.655 ;
        RECT 22.380 -10.050 22.600 -9.995 ;
        RECT 19.410 -10.250 21.500 -10.050 ;
        RECT 21.700 -10.250 22.600 -10.050 ;
        RECT 19.410 -10.435 19.640 -10.250 ;
        RECT 11.830 -10.900 15.050 -10.700 ;
        RECT 11.830 -11.065 12.525 -10.900 ;
        RECT 16.090 -11.065 16.420 -10.435 ;
        RECT 19.310 -11.065 19.640 -10.435 ;
        RECT 22.380 -10.575 22.600 -10.250 ;
        RECT 22.785 -10.725 22.965 -9.825 ;
        RECT 23.135 -10.555 23.510 -9.995 ;
        RECT 23.715 -10.065 24.025 -9.995 ;
        RECT 25.500 -10.065 26.350 -10.050 ;
        RECT 26.730 -10.065 27.060 -10.005 ;
        RECT 23.715 -10.235 24.780 -10.065 ;
        RECT 25.500 -10.235 27.060 -10.065 ;
        RECT 23.715 -10.325 24.025 -10.235 ;
        RECT 25.500 -10.250 26.350 -10.235 ;
        RECT 26.730 -10.245 27.060 -10.235 ;
        RECT 23.685 -10.725 24.015 -10.495 ;
        RECT 22.785 -10.750 24.015 -10.725 ;
        RECT 26.150 -10.750 26.350 -10.250 ;
        RECT 22.785 -10.950 26.350 -10.750 ;
        RECT 22.785 -11.065 24.015 -10.950 ;
        RECT 10.855 -12.350 11.550 -11.965 ;
        RECT 14.085 -12.200 14.780 -12.025 ;
        RECT 9.800 -12.550 11.550 -12.350 ;
        RECT 10.855 -12.595 11.550 -12.550 ;
        RECT 10.875 -12.865 11.210 -12.785 ;
        RECT 9.565 -13.035 11.210 -12.865 ;
        RECT 11.380 -13.195 11.550 -12.595 ;
        RECT 12.350 -12.400 14.780 -12.200 ;
        RECT 11.720 -12.800 12.055 -12.765 ;
        RECT 12.350 -12.800 12.550 -12.400 ;
        RECT 11.720 -13.000 12.550 -12.800 ;
        RECT 11.720 -13.035 12.055 -13.000 ;
        RECT 11.285 -14.175 11.615 -13.195 ;
        RECT 12.900 -13.700 13.100 -12.400 ;
        RECT 14.085 -12.655 14.780 -12.400 ;
        RECT 14.105 -12.865 14.440 -12.845 ;
        RECT 13.565 -13.035 14.440 -12.865 ;
        RECT 14.105 -13.095 14.440 -13.035 ;
        RECT 14.610 -13.255 14.780 -12.655 ;
        RECT 14.950 -12.850 15.285 -12.825 ;
        RECT 14.950 -13.050 16.700 -12.850 ;
        RECT 14.950 -13.095 15.285 -13.050 ;
        RECT 14.515 -14.235 14.845 -13.255 ;
      LAYER met1 ;
        RECT 12.120 6.550 12.380 6.610 ;
        RECT 24.340 6.550 24.660 6.580 ;
        RECT 12.120 6.350 24.660 6.550 ;
        RECT 12.120 6.290 12.380 6.350 ;
        RECT 24.340 6.320 24.660 6.350 ;
        RECT 12.090 3.620 12.410 3.880 ;
        RECT 24.370 3.840 24.630 4.160 ;
        RECT 19.840 3.800 20.160 3.830 ;
        RECT 12.150 2.915 12.350 3.620 ;
        RECT 13.150 3.100 13.450 3.780 ;
        RECT 19.840 3.600 22.450 3.800 ;
        RECT 19.840 3.570 20.160 3.600 ;
        RECT 12.105 2.685 12.395 2.915 ;
        RECT 13.120 2.800 13.480 3.100 ;
        RECT 22.250 2.845 22.450 3.600 ;
        RECT 24.400 3.510 24.600 3.840 ;
        RECT 24.370 3.190 24.630 3.510 ;
        RECT 22.235 2.555 22.465 2.845 ;
        RECT 23.825 2.630 24.085 2.665 ;
        RECT 23.795 2.375 24.110 2.630 ;
        RECT 23.825 2.345 24.085 2.375 ;
        RECT 19.640 2.000 19.960 2.030 ;
        RECT 20.705 2.000 20.995 2.015 ;
        RECT 19.640 1.800 20.995 2.000 ;
        RECT 19.640 1.770 19.960 1.800 ;
        RECT 20.705 1.785 20.995 1.800 ;
        RECT 11.520 -0.010 11.780 0.310 ;
        RECT 12.120 -0.010 12.380 0.310 ;
        RECT 14.940 0.170 15.260 0.430 ;
        RECT 12.150 -0.390 12.350 -0.010 ;
        RECT 8.355 -0.665 8.645 -0.435 ;
        RECT 8.400 -3.550 8.600 -0.665 ;
        RECT 11.410 -0.720 11.670 -0.690 ;
        RECT 12.120 -0.710 12.380 -0.390 ;
        RECT 12.620 -0.660 12.880 -0.340 ;
        RECT 15.020 -0.355 15.180 0.170 ;
        RECT 15.670 -0.060 15.930 0.260 ;
        RECT 19.640 0.170 19.960 0.430 ;
        RECT 14.985 -0.645 15.215 -0.355 ;
        RECT 11.380 -0.980 11.670 -0.720 ;
        RECT 11.410 -1.010 11.670 -0.980 ;
        RECT 11.445 -1.655 11.765 -1.615 ;
        RECT 12.660 -1.655 12.845 -0.660 ;
        RECT 11.445 -1.840 12.845 -1.655 ;
        RECT 11.445 -1.875 11.765 -1.840 ;
        RECT 15.700 -3.550 15.900 -0.060 ;
        RECT 19.700 -0.150 19.900 0.170 ;
        RECT 19.700 -0.350 24.850 -0.150 ;
        RECT 18.570 -1.010 18.830 -0.690 ;
        RECT 18.600 -1.555 18.800 -1.010 ;
        RECT 18.585 -1.845 18.815 -1.555 ;
        RECT 19.320 -2.250 19.580 -2.190 ;
        RECT 19.320 -2.450 20.950 -2.250 ;
        RECT 19.320 -2.510 19.580 -2.450 ;
        RECT 20.750 -2.905 20.950 -2.450 ;
        RECT 24.650 -2.905 24.850 -0.350 ;
        RECT 17.605 -3.165 17.895 -2.935 ;
        RECT 8.400 -3.750 15.900 -3.550 ;
        RECT 11.450 -4.275 11.770 -4.015 ;
        RECT 11.520 -5.545 11.705 -4.275 ;
        RECT 13.640 -4.790 13.960 -4.770 ;
        RECT 17.640 -4.790 17.860 -3.165 ;
        RECT 20.735 -3.195 20.965 -2.905 ;
        RECT 24.635 -3.195 24.865 -2.905 ;
        RECT 21.710 -3.500 22.000 -3.475 ;
        RECT 22.425 -3.500 22.685 -3.435 ;
        RECT 19.570 -3.600 19.830 -3.540 ;
        RECT 21.105 -3.600 21.395 -3.585 ;
        RECT 19.570 -3.800 21.395 -3.600 ;
        RECT 21.710 -3.685 22.685 -3.500 ;
        RECT 21.710 -3.705 22.000 -3.685 ;
        RECT 22.425 -3.755 22.685 -3.685 ;
        RECT 19.570 -3.860 19.830 -3.800 ;
        RECT 21.105 -3.815 21.395 -3.800 ;
        RECT 13.640 -5.010 17.860 -4.790 ;
        RECT 18.655 -4.955 18.945 -4.935 ;
        RECT 20.640 -4.955 20.960 -4.920 ;
        RECT 13.640 -5.030 13.960 -5.010 ;
        RECT 18.655 -5.145 20.960 -4.955 ;
        RECT 18.655 -5.165 18.945 -5.145 ;
        RECT 20.640 -5.180 20.960 -5.145 ;
        RECT 23.140 -5.545 23.460 -5.505 ;
        RECT 11.520 -5.730 23.460 -5.545 ;
        RECT 11.520 -7.405 11.705 -5.730 ;
        RECT 23.140 -5.765 23.460 -5.730 ;
        RECT 5.660 -7.590 11.705 -7.405 ;
        RECT 13.050 -6.600 25.700 -6.400 ;
        RECT 13.050 -7.490 13.250 -6.600 ;
        RECT 25.500 -7.470 25.700 -6.600 ;
        RECT 5.665 -14.570 5.835 -7.590 ;
        RECT 13.020 -7.810 13.280 -7.490 ;
        RECT 25.440 -7.730 25.760 -7.470 ;
        RECT 12.990 -9.330 13.310 -9.070 ;
        RECT 21.250 -9.250 23.450 -9.050 ;
        RECT 13.050 -9.985 13.250 -9.330 ;
        RECT 14.170 -9.580 14.430 -9.260 ;
        RECT 13.640 -9.800 13.960 -9.770 ;
        RECT 14.200 -9.800 14.400 -9.580 ;
        RECT 13.005 -10.215 13.295 -9.985 ;
        RECT 13.640 -10.000 14.400 -9.800 ;
        RECT 13.640 -10.030 13.960 -10.000 ;
        RECT 14.200 -10.235 14.400 -10.000 ;
        RECT 21.250 -10.020 21.450 -9.250 ;
        RECT 14.155 -10.465 14.445 -10.235 ;
        RECT 21.190 -10.280 21.510 -10.020 ;
        RECT 21.655 -10.265 21.945 -10.035 ;
        RECT 23.250 -10.055 23.450 -9.250 ;
        RECT 24.535 -9.330 24.855 -9.070 ;
        RECT 25.470 -9.310 25.730 -8.990 ;
        RECT 24.610 -10.005 24.780 -9.330 ;
        RECT 25.500 -9.990 25.700 -9.310 ;
        RECT 21.700 -10.620 21.900 -10.265 ;
        RECT 23.235 -10.345 23.465 -10.055 ;
        RECT 24.580 -10.295 24.810 -10.005 ;
        RECT 25.470 -10.310 25.730 -9.990 ;
        RECT 21.640 -10.880 21.960 -10.620 ;
        RECT 9.770 -12.610 10.030 -12.290 ;
        RECT 13.490 -12.480 13.810 -12.220 ;
        RECT 16.470 -12.410 16.730 -12.090 ;
        RECT 13.565 -12.805 13.735 -12.480 ;
        RECT 9.505 -13.065 9.795 -12.835 ;
        RECT 9.570 -14.570 9.730 -13.065 ;
        RECT 13.535 -13.095 13.765 -12.805 ;
        RECT 16.500 -12.820 16.700 -12.410 ;
        RECT 20.670 -12.460 20.930 -12.140 ;
        RECT 16.440 -13.080 16.760 -12.820 ;
        RECT 12.840 -13.500 13.160 -13.470 ;
        RECT 20.700 -13.500 20.900 -12.460 ;
        RECT 21.670 -12.560 21.930 -12.240 ;
        RECT 21.700 -13.500 21.900 -12.560 ;
        RECT 12.840 -13.700 21.900 -13.500 ;
        RECT 12.840 -13.730 13.160 -13.700 ;
        RECT 5.665 -14.730 9.730 -14.570 ;
        RECT 5.665 -14.735 5.835 -14.730 ;
      LAYER met2 ;
        RECT 12.090 6.320 12.410 6.580 ;
        RECT 12.150 3.910 12.350 6.320 ;
        RECT 24.370 6.290 24.630 6.610 ;
        RECT 24.400 4.130 24.600 6.290 ;
        RECT 12.120 3.590 12.380 3.910 ;
        RECT 24.340 3.870 24.660 4.130 ;
        RECT 12.110 1.850 12.390 1.885 ;
        RECT 13.150 1.850 13.450 3.130 ;
        RECT 23.795 2.375 24.115 2.635 ;
        RECT 12.100 1.550 13.450 1.850 ;
        RECT 19.670 1.740 19.930 2.060 ;
        RECT 12.110 1.515 12.390 1.550 ;
        RECT 19.700 1.200 19.900 1.740 ;
        RECT 11.550 1.000 19.900 1.200 ;
        RECT 11.550 0.280 11.750 1.000 ;
        RECT 15.000 0.460 15.200 1.000 ;
        RECT 19.700 0.460 19.900 1.000 ;
        RECT 12.100 0.280 12.400 0.345 ;
        RECT 11.490 0.020 11.810 0.280 ;
        RECT 12.090 0.020 12.410 0.280 ;
        RECT 14.970 0.140 15.230 0.460 ;
        RECT 19.670 0.140 19.930 0.460 ;
        RECT 12.100 -0.045 12.400 0.020 ;
        RECT 23.860 -0.495 24.055 2.375 ;
        RECT 11.380 -0.750 11.700 -0.720 ;
        RECT 18.540 -0.750 18.860 -0.720 ;
        RECT 11.380 -0.950 18.860 -0.750 ;
        RECT 11.380 -0.980 11.700 -0.950 ;
        RECT 18.540 -0.980 18.860 -0.950 ;
        RECT 11.475 -1.905 11.735 -1.585 ;
        RECT 11.515 -3.985 11.700 -1.905 ;
        RECT 22.395 -3.505 22.715 -3.465 ;
        RECT 23.865 -3.505 24.050 -0.495 ;
        RECT 22.395 -3.690 24.050 -3.505 ;
        RECT 22.395 -3.725 22.715 -3.690 ;
        RECT 11.480 -4.305 11.740 -3.985 ;
        RECT 13.670 -5.060 13.930 -4.740 ;
        RECT 13.690 -7.360 13.910 -5.060 ;
        RECT 20.670 -5.210 20.930 -4.890 ;
        RECT 12.990 -7.780 13.310 -7.520 ;
        RECT 13.050 -9.040 13.250 -7.780 ;
        RECT 13.020 -9.360 13.280 -9.040 ;
        RECT 13.700 -9.740 13.900 -7.360 ;
        RECT 14.140 -9.320 14.460 -9.290 ;
        RECT 14.760 -9.320 16.700 -9.300 ;
        RECT 14.140 -9.500 16.700 -9.320 ;
        RECT 14.140 -9.520 14.910 -9.500 ;
        RECT 14.140 -9.550 14.460 -9.520 ;
        RECT 13.670 -10.060 13.930 -9.740 ;
        RECT 9.800 -11.500 13.750 -11.300 ;
        RECT 9.800 -12.320 10.000 -11.500 ;
        RECT 13.550 -12.190 13.750 -11.500 ;
        RECT 16.500 -12.120 16.700 -9.500 ;
        RECT 9.740 -12.580 10.060 -12.320 ;
        RECT 13.520 -12.510 13.780 -12.190 ;
        RECT 16.440 -12.380 16.760 -12.120 ;
        RECT 20.700 -12.170 20.900 -5.210 ;
        RECT 23.170 -5.540 23.430 -5.475 ;
        RECT 23.865 -5.540 24.050 -3.690 ;
        RECT 23.170 -5.725 24.050 -5.540 ;
        RECT 23.170 -5.795 23.430 -5.725 ;
        RECT 23.865 -7.305 24.050 -5.725 ;
        RECT 23.865 -7.490 24.790 -7.305 ;
        RECT 24.610 -9.040 24.780 -7.490 ;
        RECT 25.470 -7.760 25.730 -7.440 ;
        RECT 25.500 -9.020 25.700 -7.760 ;
        RECT 24.565 -9.360 24.825 -9.040 ;
        RECT 25.440 -9.280 25.760 -9.020 ;
        RECT 21.670 -10.910 21.930 -10.590 ;
        RECT 20.640 -12.430 20.960 -12.170 ;
        RECT 21.700 -12.270 21.900 -10.910 ;
        RECT 21.640 -12.530 21.960 -12.270 ;
      LAYER met3 ;
        RECT 12.085 1.535 12.415 1.865 ;
        RECT 12.100 0.325 12.400 1.535 ;
        RECT 12.075 -0.025 12.425 0.325 ;
  END
END pfd_lay
END LIBRARY

