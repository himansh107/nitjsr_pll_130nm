magic
tech sky130A
magscale 1 2
timestamp 1714832304
<< dnwell >>
rect 1600 3810 2602 4736
rect 6342 2116 7344 3042
rect 1812 894 2814 1820
rect 4076 1156 5078 2082
<< nwell >>
rect 1882 4818 2310 5148
rect 1870 4816 2310 4818
rect 1520 4530 2682 4816
rect 1520 4016 1806 4530
rect 2396 4016 2682 4530
rect 1520 3730 2682 4016
rect 6262 2836 7424 3122
rect 2060 1900 2488 2776
rect 6262 2322 6548 2836
rect 7138 2322 7424 2836
rect 1732 1614 2894 1900
rect 1732 1100 2018 1614
rect 2608 1100 2894 1614
rect 1732 814 2894 1100
rect 3996 1876 5158 2162
rect 6262 2036 7424 2322
rect 3996 1362 4282 1876
rect 4872 1362 5158 1876
rect 3996 1076 5158 1362
<< nsubdiff >>
rect 1557 4759 2645 4779
rect 1557 4725 1637 4759
rect 2565 4725 2645 4759
rect 1557 4705 2645 4725
rect 1557 4699 1631 4705
rect 1557 3847 1577 4699
rect 1611 3847 1631 4699
rect 1557 3841 1631 3847
rect 2571 4699 2645 4705
rect 2571 3847 2591 4699
rect 2625 3847 2645 4699
rect 2571 3841 2645 3847
rect 1557 3821 2645 3841
rect 1557 3787 1637 3821
rect 2565 3787 2645 3821
rect 1557 3767 2645 3787
rect 6299 3065 7387 3085
rect 6299 3031 6379 3065
rect 7307 3031 7387 3065
rect 6299 3011 7387 3031
rect 6299 3005 6373 3011
rect 6299 2153 6319 3005
rect 6353 2153 6373 3005
rect 6299 2147 6373 2153
rect 7313 3005 7387 3011
rect 7313 2153 7333 3005
rect 7367 2153 7387 3005
rect 7313 2147 7387 2153
rect 6299 2127 7387 2147
rect 4033 2105 5121 2125
rect 4033 2071 4113 2105
rect 5041 2071 5121 2105
rect 6299 2093 6379 2127
rect 7307 2093 7387 2127
rect 6299 2073 7387 2093
rect 4033 2051 5121 2071
rect 4033 2045 4107 2051
rect 1769 1843 2857 1863
rect 1769 1809 1849 1843
rect 2777 1809 2857 1843
rect 1769 1789 2857 1809
rect 1769 1783 1843 1789
rect 1769 931 1789 1783
rect 1823 931 1843 1783
rect 1769 925 1843 931
rect 2783 1783 2857 1789
rect 2783 931 2803 1783
rect 2837 931 2857 1783
rect 4033 1193 4053 2045
rect 4087 1193 4107 2045
rect 4033 1187 4107 1193
rect 5047 2045 5121 2051
rect 5047 1193 5067 2045
rect 5101 1193 5121 2045
rect 5047 1187 5121 1193
rect 4033 1167 5121 1187
rect 4033 1133 4113 1167
rect 5041 1133 5121 1167
rect 4033 1113 5121 1133
rect 2783 925 2857 931
rect 1769 905 2857 925
rect 1769 871 1849 905
rect 2777 871 2857 905
rect 1769 851 2857 871
<< nsubdiffcont >>
rect 1637 4725 2565 4759
rect 1577 3847 1611 4699
rect 2591 3847 2625 4699
rect 1637 3787 2565 3821
rect 6379 3031 7307 3065
rect 6319 2153 6353 3005
rect 7333 2153 7367 3005
rect 4113 2071 5041 2105
rect 6379 2093 7307 2127
rect 1849 1809 2777 1843
rect 1789 931 1823 1783
rect 2803 931 2837 1783
rect 4053 1193 4087 2045
rect 5067 1193 5101 2045
rect 4113 1133 5041 1167
rect 1849 871 2777 905
<< locali >>
rect 1577 4725 1637 4759
rect 2565 4725 2625 4759
rect 1577 4699 1611 4725
rect 1577 3821 1611 3847
rect 2591 4699 2625 4725
rect 2591 3821 2625 3847
rect 1577 3787 1637 3821
rect 2565 3787 2625 3821
rect 6319 3031 6379 3065
rect 7307 3031 7367 3065
rect 6319 3005 6353 3031
rect 6319 2127 6353 2153
rect 7333 3005 7367 3031
rect 7333 2127 7367 2153
rect 4053 2071 4113 2105
rect 5041 2071 5101 2105
rect 6319 2093 6379 2127
rect 7307 2093 7367 2127
rect 4053 2045 4087 2071
rect 1789 1809 1849 1843
rect 2777 1809 2837 1843
rect 1789 1783 1823 1809
rect 1789 905 1823 931
rect 2803 1783 2837 1809
rect 4053 1167 4087 1193
rect 5067 2045 5101 2071
rect 5067 1167 5101 1193
rect 4053 1133 4113 1167
rect 5041 1133 5101 1167
rect 2803 905 2837 931
rect 1789 871 1849 905
rect 2777 871 2837 905
<< metal1 >>
rect 14936 19604 16996 19692
rect 17084 19604 17090 19692
rect 13728 17436 14580 17540
rect 14684 17436 14690 17540
rect 13728 14580 13832 17436
rect 13722 14380 14464 14580
rect 14664 14380 14670 14580
rect 13728 13352 13832 14380
rect 13722 13248 13728 13352
rect 13832 13248 13838 13352
rect 12310 12782 12414 12788
rect 12414 12678 14554 12782
rect 12310 12672 12414 12678
rect 13728 12484 13832 12490
rect 13728 9496 13832 12380
rect 12852 9392 12858 9496
rect 12962 9392 13832 9496
rect 14450 9090 14554 12678
rect 11512 8986 14554 9090
rect 11512 8746 11616 8986
rect 11520 8482 11584 8746
rect 11520 7174 11584 7502
rect 11520 7104 11580 7174
rect 11512 7016 11580 7104
rect 7824 6949 7870 6958
rect 7824 6903 8359 6949
rect -1036 6380 -980 6656
rect 7824 6652 7870 6903
rect 8313 6810 8359 6903
rect 11520 6936 11580 7016
rect 2422 6478 2474 6588
rect 2422 6420 2474 6426
rect 2774 6380 2806 6384
rect 8096 6380 8152 6650
rect 8196 6446 8398 6810
rect -1036 6324 8152 6380
rect 2416 6210 2422 6262
rect 2474 6210 2676 6262
rect 2728 6210 2734 6262
rect 1770 5944 1970 6022
rect -750 5874 1970 5944
rect 2774 5918 2806 6324
rect 2932 6262 2984 6268
rect 2984 6210 5184 6262
rect 2932 6204 2984 6210
rect 3844 6039 3910 6042
rect 3844 5973 4491 6039
rect 4557 5973 4563 6039
rect -750 3073 -680 5874
rect 1770 5800 1970 5874
rect 2758 5866 2764 5918
rect 2816 5866 2822 5918
rect 3844 5852 3910 5973
rect 3810 5800 3910 5852
rect 280 5794 3910 5800
rect 280 5690 3926 5794
rect 128 5568 134 5620
rect 186 5614 192 5620
rect 298 5614 670 5690
rect 186 5576 670 5614
rect 186 5574 380 5576
rect 186 5568 192 5574
rect 1664 5524 1720 5690
rect 3847 5669 3926 5690
rect 4332 5669 4338 5674
rect 3847 5627 4338 5669
rect 2764 5602 2816 5608
rect 2764 5544 2816 5550
rect -76 5470 506 5516
rect 1660 5472 2128 5524
rect -76 5275 -30 5470
rect 1660 5452 1720 5472
rect 128 5352 134 5404
rect 186 5398 192 5404
rect 186 5358 436 5398
rect 186 5352 192 5358
rect 500 5348 748 5392
rect -76 5229 497 5275
rect -486 5098 -286 5172
rect -76 5098 -30 5229
rect -486 5054 -30 5098
rect -486 4972 -286 5054
rect -188 3640 -144 5054
rect -76 4933 -30 5054
rect 220 5052 226 5104
rect 278 5100 284 5104
rect 704 5100 748 5348
rect 1660 5290 1712 5452
rect 1660 5232 1712 5238
rect 1818 5368 2066 5400
rect 2126 5370 2398 5412
rect 1818 5118 1850 5368
rect 1898 5290 1950 5296
rect 1950 5238 2130 5290
rect 1898 5232 1950 5238
rect 1900 5128 2278 5166
rect 1900 5118 2250 5128
rect 278 5056 1368 5100
rect 1818 5086 2250 5118
rect 2244 5076 2250 5086
rect 2302 5076 2308 5128
rect 278 5052 284 5056
rect -76 4887 505 4933
rect 1324 4896 1368 5056
rect 2356 4905 2398 5370
rect 2488 5128 2540 5134
rect 2488 5070 2540 5076
rect 1671 4896 2398 4905
rect -76 4729 -30 4887
rect 1324 4863 2398 4896
rect 2498 4936 2530 5070
rect 2774 4936 2806 5544
rect 4039 5535 4081 5627
rect 4332 5622 4338 5627
rect 4390 5622 4396 5674
rect 4739 5594 4785 6210
rect 5148 5710 5184 6210
rect 8285 6181 8351 6446
rect 6751 6115 8351 6181
rect 5307 6039 5373 6045
rect 6751 6039 6817 6115
rect 5373 5973 6817 6039
rect 5307 5967 5373 5973
rect 11520 5944 11584 6936
rect 7342 5880 11584 5944
rect 5148 5674 5322 5710
rect 5148 5636 5184 5674
rect 5140 5630 5192 5636
rect 4736 5588 4788 5594
rect 5286 5602 5322 5674
rect 5140 5572 5192 5578
rect 5260 5560 5444 5602
rect 4736 5530 4788 5536
rect 4128 5430 4508 5480
rect 4458 5365 4508 5430
rect 4910 5454 5334 5502
rect 4910 5365 4958 5454
rect 4332 5354 4338 5359
rect 2498 4904 2806 4936
rect 3868 5304 4124 5344
rect 4188 5312 4338 5354
rect 4332 5307 4338 5312
rect 4390 5307 4396 5359
rect 4458 5315 4958 5365
rect 5134 5326 5140 5378
rect 5192 5370 5198 5378
rect 5192 5334 5272 5370
rect 5351 5342 5642 5384
rect 5192 5326 5198 5334
rect 1324 4852 1713 4863
rect 220 4774 226 4826
rect 278 4822 284 4826
rect 278 4778 440 4822
rect 500 4792 754 4842
rect 278 4774 284 4778
rect -76 4683 505 4729
rect 704 4639 754 4792
rect 521 4630 754 4639
rect 302 4589 754 4630
rect 302 4496 674 4589
rect 308 3640 314 3644
rect -188 3596 314 3640
rect 308 3592 314 3596
rect 366 3592 372 3644
rect 448 3350 504 4496
rect 1540 4400 1596 4406
rect 1370 4344 1540 4400
rect 1370 4204 1426 4344
rect 1540 4338 1596 4344
rect 1671 4289 1713 4852
rect 1758 4344 1764 4400
rect 1820 4344 2136 4400
rect 1671 4247 2067 4289
rect 2498 4278 2530 4904
rect 3868 4794 3908 5304
rect 4458 5256 4508 5315
rect 4910 5264 4958 5315
rect 4458 5249 4514 5256
rect 4131 5199 4514 5249
rect 4910 5216 5328 5264
rect 4474 4794 4514 5199
rect 4736 5206 4788 5212
rect 4736 5148 4788 5154
rect 2136 4246 2530 4278
rect 2984 4754 4514 4794
rect 1370 4148 2138 4204
rect 614 3644 666 3650
rect 1176 3640 1182 3644
rect 666 3596 1182 3640
rect 1176 3592 1182 3596
rect 1234 3592 1240 3644
rect 614 3586 666 3592
rect 1370 3350 1426 4148
rect 2358 4094 2390 4246
rect 2196 4062 2390 4094
rect 2984 3814 3024 4754
rect 3204 3958 3748 4002
rect 2978 3808 3030 3814
rect 2978 3750 3030 3756
rect 3204 3754 3248 3958
rect 4739 3892 4785 5148
rect 5600 4204 5642 5342
rect 7342 4204 7406 5880
rect 14936 4824 15024 19604
rect 15562 14580 15762 14586
rect 15562 14374 15762 14380
rect 8106 4736 15024 4824
rect 8106 4204 8194 4736
rect 15618 4452 15706 14374
rect 9460 4364 15706 4452
rect 8992 4204 9192 4246
rect 5594 4132 9192 4204
rect 3654 3846 4785 3892
rect 3200 3710 3756 3754
rect 1546 3644 1598 3650
rect 3200 3640 3244 3710
rect 1598 3596 3244 3640
rect 1546 3586 1598 3592
rect 2972 3416 2978 3468
rect 3030 3416 3036 3468
rect 2984 3350 3024 3416
rect 442 3341 3056 3350
rect -389 3279 3056 3341
rect -756 3003 -750 3073
rect -680 3003 -674 3073
rect -389 694 -327 3279
rect 442 3246 3056 3279
rect -145 3177 -75 3183
rect 1404 3177 1604 3204
rect -75 3107 1604 3177
rect -145 3101 -75 3107
rect 1404 3002 1604 3107
rect 3219 3021 5307 3067
rect 472 2972 3044 3002
rect 448 2971 3044 2972
rect 3219 2971 3265 3021
rect 448 2968 3265 2971
rect 348 2928 3265 2968
rect 348 2854 388 2928
rect 448 2925 3265 2928
rect 448 2916 3044 2925
rect 336 2802 342 2854
rect 394 2802 400 2854
rect 448 2822 824 2916
rect 128 2710 634 2752
rect 1678 2736 1734 2916
rect 5261 2879 5307 3021
rect 4747 2833 5389 2879
rect 5048 2768 5090 2833
rect 1798 2736 2306 2768
rect 1678 2712 2306 2736
rect 4496 2724 4738 2760
rect 4796 2726 5090 2768
rect 128 2503 170 2710
rect 1678 2680 1854 2712
rect 336 2582 342 2634
rect 394 2628 400 2634
rect 394 2588 566 2628
rect 634 2590 894 2628
rect 394 2582 400 2588
rect 128 2461 639 2503
rect -248 2320 -48 2360
rect 128 2320 170 2461
rect -248 2264 170 2320
rect 856 2352 894 2590
rect 1798 2534 1854 2680
rect 1798 2472 1854 2478
rect 1968 2594 2240 2630
rect 2310 2616 2610 2650
rect 1968 2362 2004 2594
rect 2036 2534 2092 2540
rect 2092 2478 2320 2534
rect 2036 2472 2092 2478
rect 2084 2396 2452 2400
rect 2084 2370 2472 2396
rect 2084 2362 2466 2370
rect 856 2296 1680 2352
rect 1968 2326 2466 2362
rect 856 2265 894 2296
rect -248 2160 -48 2264
rect 6 948 62 2264
rect 128 2051 170 2264
rect 387 2227 894 2265
rect 387 2186 425 2227
rect 380 2180 432 2186
rect 380 2122 432 2128
rect 128 2009 619 2051
rect 1624 2049 1680 2296
rect 2454 2318 2466 2326
rect 2518 2318 2524 2370
rect 2454 2136 2490 2318
rect 2446 2130 2498 2136
rect 2446 2072 2498 2078
rect 1624 2039 2006 2049
rect 2576 2039 2610 2616
rect 4496 2554 4532 2724
rect 4876 2658 5069 2669
rect 4741 2623 5069 2658
rect 5023 2601 5069 2623
rect 5343 2601 5389 2833
rect 5600 2859 5642 4132
rect 8992 4042 9192 4132
rect 9460 3414 9548 4364
rect 7568 3326 9548 3414
rect 6558 2859 6564 2864
rect 5600 2817 6564 2859
rect 6558 2812 6564 2817
rect 6616 2812 6622 2864
rect 5938 2658 6892 2704
rect 5938 2601 5984 2658
rect 5023 2555 5984 2601
rect 3426 2518 4674 2554
rect 3426 2462 3462 2518
rect 5938 2499 5984 2555
rect 6558 2554 6564 2606
rect 6616 2601 6622 2606
rect 6616 2559 6819 2601
rect 6881 2575 7107 2613
rect 6616 2554 6622 2559
rect 3418 2456 3470 2462
rect 5938 2453 6891 2499
rect 3418 2398 3470 2404
rect 7069 2397 7107 2575
rect 2656 2370 2708 2376
rect 2708 2326 3846 2362
rect 2656 2312 2708 2318
rect 3412 2192 3418 2244
rect 3470 2192 3476 2244
rect 1624 2016 2610 2039
rect 128 1853 170 2009
rect 1624 2004 1680 2016
rect 1917 2005 2610 2016
rect 374 1916 380 1968
rect 432 1961 438 1968
rect 432 1923 547 1961
rect 432 1916 438 1923
rect 602 1920 850 1962
rect 128 1811 605 1853
rect 808 1767 850 1920
rect 647 1764 850 1767
rect 408 1725 850 1764
rect 408 1620 758 1725
rect 6 892 464 948
rect 520 892 526 948
rect 578 694 640 1620
rect 1810 1481 1862 1487
rect 1639 1430 1810 1480
rect 1639 1370 1689 1430
rect 1810 1423 1862 1429
rect 1486 1320 1690 1370
rect 1917 1355 1951 2005
rect 2440 1884 2446 1936
rect 2498 1884 2504 1936
rect 2020 1429 2026 1481
rect 2078 1480 2084 1481
rect 2078 1430 2328 1480
rect 2078 1429 2084 1430
rect 2454 1362 2490 1884
rect 1917 1321 2257 1355
rect 2336 1326 2490 1362
rect 740 948 795 954
rect 795 893 1378 948
rect 1433 893 1439 948
rect 740 887 795 893
rect 1486 694 1536 1320
rect 1639 1269 1689 1320
rect 2454 1288 2490 1326
rect 1639 1219 2331 1269
rect 2386 1252 2490 1288
rect 2386 1134 2422 1252
rect 3426 1076 3462 2192
rect 3810 1622 3846 2326
rect 6943 2359 7107 2397
rect 4414 1702 4620 1738
rect 4414 1622 4450 1702
rect 3810 1586 4450 1622
rect 4512 1600 5246 1638
rect 4386 1536 4422 1586
rect 4386 1500 4616 1536
rect 5208 1123 5246 1600
rect 6943 1123 6981 2359
rect 5208 1085 6981 1123
rect 3412 1024 3418 1076
rect 3470 1024 3476 1076
rect 1596 948 1651 954
rect 1651 893 3767 948
rect 1596 887 1651 893
rect 3412 768 3418 820
rect 3470 768 3476 820
rect -389 684 3386 694
rect 3426 684 3462 768
rect -389 634 3488 684
rect -389 632 1794 634
rect 2218 632 3488 634
rect 1366 -950 1454 632
rect 2721 168 2783 632
rect 2916 333 2954 340
rect 3712 333 3767 893
rect 5208 490 5246 1085
rect 5201 484 5253 490
rect 5201 426 5253 432
rect 2916 295 6053 333
rect 2721 99 2856 168
rect 2740 -160 2856 99
rect 2916 -26 2954 295
rect 3712 283 3767 295
rect 5195 192 5201 244
rect 5253 192 5259 244
rect 5208 43 5246 192
rect 2802 -232 2842 -160
rect 3056 -232 3096 -6
rect 6015 -7 6053 295
rect 2802 -272 3096 -232
rect 1366 -956 7498 -950
rect 7568 -956 7656 3326
rect 1366 -1038 7656 -956
rect 7064 -1044 7656 -1038
<< via1 >>
rect 16996 19604 17084 19692
rect 14580 17436 14684 17540
rect 14464 14380 14664 14580
rect 13728 13248 13832 13352
rect 12310 12678 12414 12782
rect 13728 12380 13832 12484
rect 12858 9392 12962 9496
rect 2422 6426 2474 6478
rect 2422 6210 2474 6262
rect 2676 6210 2728 6262
rect 2932 6210 2984 6262
rect 4491 5973 4557 6039
rect 2764 5866 2816 5918
rect 134 5568 186 5620
rect 2764 5550 2816 5602
rect 134 5352 186 5404
rect 226 5052 278 5104
rect 1660 5238 1712 5290
rect 1898 5238 1950 5290
rect 2250 5076 2302 5128
rect 2488 5076 2540 5128
rect 4338 5622 4390 5674
rect 5307 5973 5373 6039
rect 4736 5536 4788 5588
rect 5140 5578 5192 5630
rect 4338 5307 4390 5359
rect 5140 5326 5192 5378
rect 226 4774 278 4826
rect 314 3592 366 3644
rect 1540 4344 1596 4400
rect 1764 4344 1820 4400
rect 4736 5154 4788 5206
rect 614 3592 666 3644
rect 1182 3592 1234 3644
rect 2978 3756 3030 3808
rect 15562 14380 15762 14580
rect 1546 3592 1598 3644
rect 2978 3416 3030 3468
rect -750 3003 -680 3073
rect -145 3107 -75 3177
rect 342 2802 394 2854
rect 342 2582 394 2634
rect 1798 2478 1854 2534
rect 2036 2478 2092 2534
rect 380 2128 432 2180
rect 2466 2318 2518 2370
rect 2446 2078 2498 2130
rect 6564 2812 6616 2864
rect 6564 2554 6616 2606
rect 3418 2404 3470 2456
rect 2656 2318 2708 2370
rect 3418 2192 3470 2244
rect 380 1916 432 1968
rect 464 892 520 948
rect 1810 1429 1862 1481
rect 2446 1884 2498 1936
rect 2026 1429 2078 1481
rect 740 893 795 948
rect 1378 893 1433 948
rect 3418 1024 3470 1076
rect 1596 893 1651 948
rect 3418 768 3470 820
rect 5201 432 5253 484
rect 5201 192 5253 244
<< metal2 >>
rect 16996 19692 17084 19698
rect 17084 19604 17322 19692
rect 17410 19604 17419 19692
rect 16996 19598 17084 19604
rect 14580 17540 14684 17546
rect 14684 17436 15428 17540
rect 15532 17436 15541 17540
rect 14580 17430 14684 17436
rect 14464 14580 14664 14586
rect 14664 14380 15562 14580
rect 15762 14380 15768 14580
rect 14464 14374 14664 14380
rect 13728 13352 13832 13358
rect 11885 12782 11979 12786
rect 11880 12777 12310 12782
rect 11880 12683 11885 12777
rect 11979 12683 12310 12777
rect 11880 12678 12310 12683
rect 12414 12678 12420 12782
rect 11885 12674 11979 12678
rect 13728 12484 13832 13248
rect 13722 12380 13728 12484
rect 13832 12380 13838 12484
rect 12858 9496 12962 9502
rect 12473 9392 12482 9496
rect 12586 9392 12858 9496
rect 12858 9386 12962 9392
rect 2416 6426 2422 6478
rect 2474 6426 2480 6478
rect 2422 6262 2474 6426
rect 2422 6204 2474 6210
rect 2676 6262 2728 6268
rect 2728 6210 2932 6262
rect 2984 6210 2990 6262
rect 2676 6204 2728 6210
rect 4491 6039 4557 6045
rect 4557 5973 5307 6039
rect 5373 5973 5379 6039
rect 4491 5967 4557 5973
rect 2764 5918 2816 5924
rect 2764 5860 2816 5866
rect 134 5620 186 5626
rect 2774 5602 2806 5860
rect 4338 5674 4390 5680
rect 4338 5616 4390 5622
rect 134 5562 186 5568
rect 140 5410 180 5562
rect 2758 5550 2764 5602
rect 2816 5550 2822 5602
rect 134 5404 186 5410
rect 4343 5365 4385 5616
rect 4730 5536 4736 5588
rect 4788 5536 4794 5588
rect 5134 5578 5140 5630
rect 5192 5578 5198 5630
rect 134 5346 186 5352
rect 4338 5359 4390 5365
rect 4338 5301 4390 5307
rect 1654 5238 1660 5290
rect 1712 5238 1898 5290
rect 1950 5238 1956 5290
rect 4739 5206 4785 5536
rect 5148 5384 5184 5578
rect 5140 5378 5192 5384
rect 5140 5320 5192 5326
rect 4730 5154 4736 5206
rect 4788 5154 4794 5206
rect 2250 5128 2302 5134
rect 226 5104 278 5110
rect 2482 5118 2488 5128
rect 2302 5086 2488 5118
rect 2482 5076 2488 5086
rect 2540 5076 2546 5128
rect 2250 5070 2302 5076
rect 226 5046 278 5052
rect 230 4832 274 5046
rect 226 4826 278 4832
rect 226 4768 278 4774
rect 1764 4400 1820 4406
rect 1534 4344 1540 4400
rect 1596 4344 1764 4400
rect 1764 4338 1820 4344
rect 2972 3756 2978 3808
rect 3030 3756 3036 3808
rect 314 3644 366 3650
rect 1182 3644 1234 3650
rect 608 3640 614 3644
rect 366 3596 614 3640
rect 608 3592 614 3596
rect 666 3592 672 3644
rect 1540 3640 1546 3644
rect 1234 3596 1546 3640
rect 1540 3592 1546 3596
rect 1598 3592 1604 3644
rect 314 3586 366 3592
rect 1182 3586 1234 3592
rect 2984 3474 3024 3756
rect 2978 3468 3030 3474
rect 2978 3410 3030 3416
rect -151 3107 -145 3177
rect -75 3107 -69 3177
rect -750 3073 -680 3079
rect -145 3073 -75 3107
rect -680 3003 -75 3073
rect -750 2997 -680 3003
rect 6564 2864 6616 2870
rect 342 2854 394 2860
rect 6564 2806 6616 2812
rect 342 2796 394 2802
rect 348 2640 388 2796
rect 342 2634 394 2640
rect 6569 2612 6611 2806
rect 342 2576 394 2582
rect 6564 2606 6616 2612
rect 6564 2548 6616 2554
rect 1792 2478 1798 2534
rect 1854 2478 2036 2534
rect 2092 2478 2098 2534
rect 3412 2404 3418 2456
rect 3470 2404 3476 2456
rect 2466 2370 2518 2376
rect 2650 2362 2656 2370
rect 2518 2326 2656 2362
rect 2650 2318 2656 2326
rect 2708 2318 2714 2370
rect 2466 2312 2518 2318
rect 3426 2250 3462 2404
rect 3418 2244 3470 2250
rect 3418 2186 3470 2192
rect 374 2128 380 2180
rect 432 2128 438 2180
rect 387 1974 425 2128
rect 2440 2078 2446 2130
rect 2498 2078 2504 2130
rect 380 1968 432 1974
rect 2454 1942 2490 2078
rect 380 1910 432 1916
rect 2446 1936 2498 1942
rect 2446 1878 2498 1884
rect 2026 1481 2078 1487
rect 1804 1429 1810 1481
rect 1862 1480 1868 1481
rect 1862 1430 2026 1480
rect 1862 1429 1868 1430
rect 2026 1423 2078 1429
rect 3418 1076 3470 1082
rect 3418 1018 3470 1024
rect 464 948 520 954
rect 1378 948 1433 954
rect 520 893 740 948
rect 795 893 801 948
rect 1433 893 1596 948
rect 1651 893 1657 948
rect 464 886 520 892
rect 1378 887 1433 893
rect 3426 826 3462 1018
rect 3418 820 3470 826
rect 3418 762 3470 768
rect 5195 432 5201 484
rect 5253 432 5259 484
rect 5208 250 5246 432
rect 5201 244 5253 250
rect 5201 186 5253 192
<< via2 >>
rect 17322 19604 17410 19692
rect 15428 17436 15532 17540
rect 11885 12683 11979 12777
rect 12482 9392 12586 9496
<< metal3 >>
rect -64956 79144 -64852 79150
rect -64956 78557 -64852 79040
rect -64961 78455 -64955 78557
rect -64853 78455 -64847 78557
rect -64956 78454 -64852 78455
rect 11360 72550 11464 72556
rect 11360 71945 11464 72446
rect 11360 71843 11361 71945
rect 11463 71843 11464 71945
rect 11360 71842 11464 71843
rect 11361 71837 11463 71842
rect -64782 65850 -64678 65856
rect -64782 65401 -64678 65746
rect -64787 65299 -64781 65401
rect -64679 65299 -64673 65401
rect -64782 65298 -64678 65299
rect 11370 59446 11474 59452
rect 11370 58785 11474 59342
rect 11365 58683 11371 58785
rect 11473 58683 11479 58785
rect 11370 58682 11474 58683
rect -64812 52654 -64708 52660
rect -64812 52175 -64708 52550
rect -64817 52073 -64811 52175
rect -64709 52073 -64703 52175
rect -64812 52072 -64708 52073
rect 11378 46084 11482 46090
rect 11378 45537 11482 45980
rect 11373 45435 11379 45537
rect 11481 45435 11487 45537
rect 11378 45434 11482 45435
rect 18551 42864 19212 42865
rect 18546 42759 18552 42864
rect 18657 42759 19212 42864
rect 18551 42758 19212 42759
rect 19319 42758 19325 42865
rect -64892 39470 -64788 39476
rect -64892 38961 -64788 39366
rect -64892 38859 -64891 38961
rect -64789 38859 -64788 38961
rect -64892 38858 -64788 38859
rect -64891 38853 -64789 38858
rect 51198 36600 51204 36704
rect 51308 36600 51314 36704
rect 51204 35839 51308 36600
rect 51199 35737 51205 35839
rect 51307 35737 51313 35839
rect 51204 35736 51308 35737
rect 11416 32862 11520 32868
rect 11416 32353 11520 32758
rect 11411 32251 11417 32353
rect 11519 32251 11525 32353
rect 11416 32250 11520 32251
rect 19128 26610 19232 26616
rect -64848 26244 -64744 26250
rect -64848 25747 -64744 26140
rect 19128 25995 19232 26506
rect 19123 25893 19129 25995
rect 19231 25893 19237 25995
rect 19128 25892 19232 25893
rect -64853 25645 -64847 25747
rect -64745 25645 -64739 25747
rect -64848 25644 -64744 25645
rect 51120 22928 51126 23032
rect 51230 23031 51762 23032
rect 51230 22929 51659 23031
rect 51761 22929 51767 23031
rect 51230 22928 51762 22929
rect 17317 19692 17415 19697
rect 11424 19604 11528 19610
rect 17317 19604 17322 19692
rect 17410 19604 17684 19692
rect 17772 19604 17778 19692
rect 17317 19599 17415 19604
rect 11424 19139 11528 19500
rect 11419 19037 11425 19139
rect 11527 19037 11533 19139
rect 11424 19036 11528 19037
rect 15423 17540 15537 17545
rect 15423 17436 15428 17540
rect 15532 17436 16584 17540
rect 16688 17436 16694 17540
rect 15423 17431 15537 17436
rect -65022 13194 -64918 13200
rect -65022 12479 -64918 13090
rect 11429 12782 11531 12787
rect 11428 12781 11984 12782
rect 11428 12679 11429 12781
rect 11531 12777 11984 12781
rect 11531 12683 11885 12777
rect 11979 12683 11984 12777
rect 11531 12679 11984 12683
rect 11428 12678 11984 12679
rect 11429 12673 11531 12678
rect -65027 12377 -65021 12479
rect -64919 12377 -64913 12479
rect -65022 12376 -64918 12377
rect 12477 9496 12591 9501
rect 11978 9392 11984 9496
rect 12088 9392 12482 9496
rect 12586 9392 12591 9496
rect 12477 9387 12591 9392
<< via3 >>
rect -64956 79040 -64852 79144
rect -64955 78455 -64853 78557
rect 11360 72446 11464 72550
rect 11361 71843 11463 71945
rect -64782 65746 -64678 65850
rect -64781 65299 -64679 65401
rect 11370 59342 11474 59446
rect 11371 58683 11473 58785
rect -64812 52550 -64708 52654
rect -64811 52073 -64709 52175
rect 11378 45980 11482 46084
rect 11379 45435 11481 45537
rect 18552 42759 18657 42864
rect 19212 42758 19319 42865
rect -64892 39366 -64788 39470
rect -64891 38859 -64789 38961
rect 51204 36600 51308 36704
rect 51205 35737 51307 35839
rect 11416 32758 11520 32862
rect 11417 32251 11519 32353
rect 19128 26506 19232 26610
rect -64848 26140 -64744 26244
rect 19129 25893 19231 25995
rect -64847 25645 -64745 25747
rect 51126 22928 51230 23032
rect 51659 22929 51761 23031
rect 11424 19500 11528 19604
rect 17684 19604 17772 19692
rect 11425 19037 11527 19139
rect 16584 17436 16688 17540
rect -65022 13090 -64918 13194
rect 11429 12679 11531 12781
rect -65021 12377 -64919 12479
rect 11984 9392 12088 9496
<< metal4 >>
rect -65492 85422 -64458 85526
rect -65492 78902 -65388 85422
rect -64956 82118 -64476 82222
rect -64956 79145 -64852 82118
rect -64957 79144 -64851 79145
rect -64957 79040 -64956 79144
rect -64852 79040 -64851 79144
rect -64957 79039 -64851 79040
rect -65492 78798 -64460 78902
rect 11184 78794 11982 78898
rect -64956 78557 -64852 78558
rect -64956 78455 -64955 78557
rect -64853 78455 -64852 78557
rect -64956 75622 -64852 78455
rect -64956 75518 -64460 75622
rect 11183 75511 11465 75617
rect 11359 72550 11465 75511
rect 11359 72446 11360 72550
rect 11464 72446 11465 72550
rect 11359 72445 11465 72446
rect 11878 72290 11982 78794
rect -65204 72176 -64450 72280
rect 11172 72186 11982 72290
rect -65204 65678 -65100 72176
rect 11360 71945 11464 71946
rect 11360 71843 11361 71945
rect 11463 71843 11464 71945
rect 11360 69010 11464 71843
rect -64782 68898 -64446 69002
rect 11172 68906 11464 69010
rect -64782 65851 -64678 68898
rect -64783 65850 -64677 65851
rect -64783 65746 -64782 65850
rect -64678 65746 -64677 65850
rect -64783 65745 -64677 65746
rect -65204 65574 -64460 65678
rect 11206 65566 12244 65670
rect -64782 65401 -64678 65402
rect -64782 65299 -64781 65401
rect -64679 65299 -64678 65401
rect -64782 62398 -64678 65299
rect -64782 62294 -64460 62398
rect 11162 62304 11474 62408
rect 11370 59447 11474 62304
rect 11369 59446 11475 59447
rect 11369 59342 11370 59446
rect 11474 59342 11475 59446
rect 11369 59341 11475 59342
rect -65058 58980 -64450 59084
rect 12140 59066 12244 65566
rect -65058 52454 -64954 58980
rect 11172 58962 12244 59066
rect 11370 58785 11474 58786
rect 11370 58683 11371 58785
rect 11473 58683 11474 58785
rect 11370 55786 11474 58683
rect -64812 55662 -64482 55766
rect 11166 55682 11474 55786
rect -64812 52655 -64708 55662
rect -64813 52654 -64707 52655
rect -64813 52550 -64812 52654
rect -64708 52550 -64707 52654
rect -64813 52549 -64707 52550
rect -65058 52350 -64460 52454
rect 11174 52358 12096 52462
rect -64812 52175 -64708 52176
rect -64812 52073 -64811 52175
rect -64709 52073 -64708 52175
rect -64812 49174 -64708 52073
rect -64812 49070 -64450 49174
rect 11208 49078 11482 49182
rect 11378 46085 11482 49078
rect 11377 46084 11483 46085
rect 11377 45980 11378 46084
rect 11482 45980 11483 46084
rect 11377 45979 11483 45980
rect 11992 45842 12096 52358
rect -65526 45738 -64476 45842
rect 11172 45738 12096 45842
rect 19020 46038 19710 46142
rect -65526 39230 -65422 45738
rect 11378 45537 11482 45538
rect 11378 45435 11379 45537
rect 11481 45435 11482 45537
rect -64892 42464 -64380 42568
rect 11378 42562 11482 45435
rect -64892 39471 -64788 42464
rect 11158 42458 11482 42562
rect 18551 42864 18658 42865
rect 18551 42759 18552 42864
rect 18657 42759 18658 42864
rect -64893 39470 -64787 39471
rect -64893 39366 -64892 39470
rect -64788 39366 -64787 39470
rect -64893 39365 -64787 39366
rect -65526 39126 -64460 39230
rect 11182 39128 11786 39232
rect -64892 38961 -64788 38962
rect -64892 38859 -64891 38961
rect -64789 38859 -64788 38961
rect -64892 35950 -64788 38859
rect -64892 35846 -64460 35950
rect 11234 35834 11520 35938
rect 11416 32863 11520 35834
rect 11415 32862 11521 32863
rect 11415 32758 11416 32862
rect 11520 32758 11521 32862
rect 11415 32757 11521 32758
rect 11682 32618 11786 39128
rect 18551 36252 18658 42759
rect 19020 39532 19124 46038
rect 19211 42865 19320 42866
rect 19211 42758 19212 42865
rect 19319 42758 19539 42865
rect 19211 42757 19320 42758
rect 19020 39428 19550 39532
rect 50964 39432 51308 39536
rect 51204 36705 51308 39432
rect 51203 36704 51309 36705
rect 51203 36600 51204 36704
rect 51308 36600 51309 36704
rect 51203 36599 51309 36600
rect 18551 36148 19550 36252
rect 50987 36150 51688 36253
rect 18551 36147 18658 36148
rect 51204 35839 51308 35840
rect 51204 35737 51205 35839
rect 51307 35737 51308 35839
rect 51204 32920 51308 35737
rect -65230 32502 -64454 32606
rect 11172 32514 11786 32618
rect 18700 32814 19554 32918
rect 50942 32816 51308 32920
rect -65230 26006 -65126 32502
rect 11416 32353 11520 32354
rect 11416 32251 11417 32353
rect 11519 32251 11520 32353
rect -64848 29240 -64480 29344
rect 11416 29338 11520 32251
rect -64848 26245 -64744 29240
rect 11172 29234 11520 29338
rect 18700 26308 18804 32814
rect 51585 29640 51688 36150
rect 19128 29526 19512 29630
rect 50942 29536 51688 29640
rect 19128 26611 19232 29526
rect 19127 26610 19233 26611
rect 19127 26506 19128 26610
rect 19232 26506 19233 26610
rect 19127 26505 19233 26506
rect -64849 26244 -64743 26245
rect -64849 26140 -64848 26244
rect -64744 26140 -64743 26244
rect 18700 26204 19550 26308
rect 51008 26216 51416 26320
rect -64849 26139 -64743 26140
rect -65230 25902 -64460 26006
rect 19128 25995 19232 25996
rect 11206 25888 11986 25992
rect -64848 25747 -64744 25748
rect -64848 25645 -64847 25747
rect -64745 25645 -64744 25747
rect -64848 22726 -64744 25645
rect -64848 22622 -64460 22726
rect 11186 22640 11528 22744
rect 11424 19605 11528 22640
rect 11423 19604 11529 19605
rect 11423 19500 11424 19604
rect 11528 19500 11529 19604
rect 11423 19499 11529 19500
rect 11882 19394 11986 25888
rect 19128 25893 19129 25995
rect 19231 25893 19232 25995
rect 19128 23028 19232 25893
rect 51125 23032 51231 23033
rect 19128 22924 19550 23028
rect 50936 22928 51126 23032
rect 51230 22928 51231 23032
rect 51125 22927 51231 22928
rect 51312 19696 51416 26216
rect 17683 19692 17773 19693
rect 17683 19604 17684 19692
rect 17772 19604 19508 19692
rect 17683 19603 17773 19604
rect 50942 19592 51416 19696
rect 51658 23031 51762 23032
rect 51658 22929 51659 23031
rect 51761 22929 51762 23031
rect -65388 19260 -64470 19364
rect 11156 19290 11986 19394
rect -65388 12782 -65284 19260
rect 11424 19139 11528 19140
rect 11424 19037 11425 19139
rect 11527 19037 11528 19139
rect -65022 16020 -64438 16124
rect 11424 16114 11528 19037
rect 16583 17540 16689 17541
rect 16583 17436 16584 17540
rect 16688 17436 19226 17540
rect 16583 17435 16689 17436
rect 19122 16412 19226 17436
rect 51658 16416 51762 22929
rect 19122 16308 19536 16412
rect 50942 16312 51762 16416
rect -65022 13195 -64918 16020
rect 11172 16010 11528 16114
rect -65023 13194 -64917 13195
rect -65023 13090 -65022 13194
rect -64918 13090 -64917 13194
rect -65023 13089 -64917 13090
rect -65388 12678 -64460 12782
rect 11172 12781 11532 12782
rect 11172 12679 11429 12781
rect 11531 12679 11532 12781
rect 11172 12678 11532 12679
rect -65022 12479 -64918 12480
rect -65022 12377 -65021 12479
rect -64919 12377 -64918 12479
rect -65022 9502 -64918 12377
rect -65022 9496 11480 9502
rect 11983 9496 12089 9497
rect -65022 9398 11984 9496
rect 11366 9392 11984 9398
rect 12088 9392 12089 9496
rect 11983 9391 12089 9392
use fd_8  fd_8_0
timestamp 1714651723
transform 1 0 14192 0 1 -282
box 2280 -462 21940 10276
use sky130_fd_pr__cap_mim_m3_1_39XMLG  sky130_fd_pr__cap_mim_m3_1_39XMLG_0
timestamp 1714629389
transform 0 1 35246 -1 0 32722
box -16410 -15800 16410 15800
use sky130_fd_pr__cap_mim_m3_1_Z926RQ  sky130_fd_pr__cap_mim_m3_1_Z926RQ_0
timestamp 1714629389
transform 0 1 -26644 -1 0 48950
box -39552 -37920 39552 37920
use sky130_fd_pr__nfet_01v8_6FB27G  sky130_fd_pr__nfet_01v8_6FB27G_0
timestamp 1714564928
transform 1 0 4588 0 1 1616
box -214 -252 214 252
use sky130_fd_pr__nfet_01v8_6FB46G  sky130_fd_pr__nfet_01v8_6FB46G_0
timestamp 1713284121
transform 1 0 474 0 1 4806
box -214 -252 214 252
use sky130_fd_pr__nfet_01v8_6FB46G  sky130_fd_pr__nfet_01v8_6FB46G_1
timestamp 1713284121
transform 1 0 6848 0 1 2582
box -214 -252 214 252
use sky130_fd_pr__nfet_01v8_6FB46G  sky130_fd_pr__nfet_01v8_6FB46G_2
timestamp 1713284121
transform 1 0 2100 0 1 4274
box -214 -252 214 252
use sky130_fd_pr__nfet_01v8_6FB46G  sky130_fd_pr__nfet_01v8_6FB46G_3
timestamp 1713284121
transform 1 0 580 0 1 1938
box -214 -252 214 252
use sky130_fd_pr__nfet_01v8_6FB46G  sky130_fd_pr__nfet_01v8_6FB46G_5
timestamp 1713284121
transform 1 0 2296 0 1 1354
box -214 -252 214 252
use sky130_fd_pr__pfet_01v8_K9S7EM  sky130_fd_pr__pfet_01v8_K9S7EM_0
timestamp 1714562015
transform 1 0 2096 0 1 5383
box -214 -273 214 273
use sky130_fd_pr__pfet_01v8_K9S7EM  sky130_fd_pr__pfet_01v8_K9S7EM_1
timestamp 1714562015
transform 1 0 2274 0 1 2627
box -214 -273 214 273
use sky130_fd_pr__pfet_01v8_KZR7FM  sky130_fd_pr__pfet_01v8_KZR7FM_0
timestamp 1714283992
transform 1 0 4158 0 1 5333
box -214 -273 214 273
use sky130_fd_pr__pfet_01v8_KZR7FM  sky130_fd_pr__pfet_01v8_KZR7FM_1
timestamp 1714283992
transform 1 0 470 0 1 5373
box -214 -273 214 273
use vco  vco_0
timestamp 1713777229
transform 1 0 7818 0 1 4469
box 442 -4993 14254 -1778
use sky130_fd_pr__nfet_01v8_HAAXKC  XM3
timestamp 1714294046
transform 0 1 4490 -1 0 12
box -214 -1710 214 1710
use sky130_fd_pr__pfet_01v8_7PMXFU  XM4
timestamp 1714283992
transform 0 1 3561 -1 0 6620
box -214 -4719 214 4719
use sky130_fd_pr__pfet_01v8_KXJ7FM  XM7
timestamp 1714283992
transform 1 0 5300 0 1 5357
box -214 -273 214 273
use sky130_fd_pr__pfet_01v8_K9S5FM  XM10
timestamp 1714285468
transform 1 0 3722 0 1 3859
box -214 -273 214 273
use sky130_fd_pr__pfet_01v8_KZR7FM  XM12
timestamp 1714283992
transform 1 0 602 0 1 2613
box -214 -273 214 273
use sky130_fd_pr__nfet_01v8_6FB46G  XM18
timestamp 1713284121
transform 1 0 4768 0 1 2738
box -214 -252 214 252
use sky130_fd_pr__res_generic_po_447X6E  XR2
timestamp 1714283992
transform 1 0 11552 0 1 7975
box -214 -761 214 761
<< labels >>
flabel metal1 -486 4972 -286 5172 0 FreeSans 256 0 0 0 up
port 0 nsew
flabel metal1 8992 4042 9192 4242 0 FreeSans 256 0 0 0 vctrl
port 1 nsew
flabel metal1 2132 662 2132 662 0 FreeSans 256 0 0 0 GND
port 10 nsew
flabel metal1 -248 2160 -48 2360 0 FreeSans 256 0 0 0 down
port 4 nsew
flabel metal1 1404 3004 1604 3204 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 1770 5822 1970 6022 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 1108 5078 1108 5078 0 FreeSans 256 0 0 0 up_bar
flabel metal1 2790 5076 2790 5076 0 FreeSans 256 0 0 0 up_bar2
flabel metal1 4760 4520 4760 4520 0 FreeSans 256 0 0 0 up_carry
flabel metal1 1154 2318 1154 2318 0 FreeSans 256 0 0 0 down_b
flabel metal1 3108 2352 3108 2352 0 FreeSans 256 0 0 0 down_b2
flabel metal1 5224 1394 5224 1394 0 FreeSans 256 0 0 0 down_carry
<< end >>
