magic
tech sky130A
magscale 1 2
timestamp 1713507270
<< nwell >>
rect 7229 986 7423 1046
<< pwell >>
rect 5002 -122 5050 8
rect 2590 -256 2762 -216
rect 3549 -610 3767 -560
rect 6136 -572 6504 -416
rect 7138 -616 7518 -490
<< viali >>
rect 3188 2542 3242 2692
rect 2474 1960 2538 2140
rect 6550 1818 6590 1994
rect -237 1012 -43 1064
rect 6228 1034 6410 1102
rect 2466 966 2654 1006
rect 3538 972 3732 1024
rect 7229 994 7423 1054
rect 1321 352 1365 522
rect 5268 420 5314 642
rect 617 -218 659 -46
rect 4582 -108 4624 86
rect 6241 -476 6407 -428
rect 2476 -526 2650 -490
rect -233 -566 -63 -526
rect 7241 -544 7413 -500
rect 3549 -610 3767 -560
<< metal1 >>
rect 2136 3865 2836 3879
rect 2136 3825 8150 3865
rect 2136 2519 2190 3825
rect 2761 3811 8150 3825
rect 2734 3010 2796 3096
rect 3069 3016 3121 3022
rect 2444 2970 3069 3010
rect 2444 2584 2484 2970
rect 2734 2968 2796 2970
rect 6754 3000 6954 3206
rect 3069 2958 3121 2964
rect 6812 2915 6876 3000
rect 2886 2860 3550 2900
rect 2886 2650 2926 2860
rect 3180 2722 3298 2784
rect 3069 2716 3121 2722
rect 3069 2662 3121 2664
rect 3180 2692 3476 2722
rect 326 2465 2190 2519
rect -253 1176 -53 1446
rect -453 1090 -447 1142
rect -395 1139 -389 1142
rect -333 1139 29 1176
rect -395 1093 29 1139
rect -395 1090 -389 1093
rect -333 1064 29 1093
rect -333 1012 -237 1064
rect -43 1012 29 1064
rect -333 1002 29 1012
rect -571 888 -105 940
rect -833 268 -633 362
rect -571 310 -519 888
rect -453 781 -447 833
rect -395 830 -389 833
rect -395 784 -173 830
rect -395 781 -389 784
rect -111 562 179 604
rect -571 268 -105 310
rect -833 258 -105 268
rect -833 210 -515 258
rect -833 156 -633 210
rect -571 -94 -519 210
rect 128 184 170 562
rect 127 126 284 184
rect 326 133 380 2465
rect 2750 2328 2786 2588
rect 3062 2576 3128 2662
rect 3180 2542 3188 2692
rect 3242 2542 3476 2692
rect 3510 2638 3550 2860
rect 6495 2857 7130 2915
rect 7188 2857 7194 2915
rect 3507 2586 4093 2638
rect 3180 2522 3476 2542
rect 3180 2494 3298 2522
rect 3510 2376 3550 2586
rect 3160 2374 3550 2376
rect 1939 2292 2786 2328
rect 3118 2336 3550 2374
rect 3118 2306 3172 2336
rect 802 934 1002 1140
rect 868 810 918 934
rect 1204 810 1256 814
rect 562 750 1258 810
rect 570 392 622 750
rect 1056 588 1108 594
rect 1056 530 1108 536
rect 1062 460 1102 530
rect 884 135 922 408
rect 1204 396 1256 750
rect 1326 706 1378 712
rect 1378 660 1694 700
rect 1326 648 1378 654
rect 1309 540 1413 574
rect 1309 522 1571 540
rect 1309 352 1321 522
rect 1365 352 1571 522
rect 1309 336 1571 352
rect 1309 260 1413 336
rect 433 133 923 135
rect -367 36 -361 88
rect -309 83 -303 88
rect 128 83 170 126
rect -309 41 170 83
rect 326 82 923 133
rect 1654 128 1694 660
rect 1939 128 1975 2292
rect 2402 2158 2550 2208
rect 2244 2140 2550 2158
rect 2244 1960 2474 2140
rect 2538 1960 2550 2140
rect 2244 1958 2550 1960
rect 2402 1890 2550 1958
rect 2602 1798 2650 2078
rect 2750 2072 2786 2292
rect 2916 2044 2968 2086
rect 2770 1942 2810 2014
rect 2916 1986 2968 1992
rect 3122 1942 3162 2306
rect 2770 1902 3162 1942
rect 2910 1798 2916 1800
rect 2602 1750 2916 1798
rect 2658 1484 2858 1750
rect 2910 1748 2916 1750
rect 2968 1748 2974 1800
rect 2462 1138 2662 1346
rect 3542 1138 3742 1384
rect 2292 1038 2298 1090
rect 2350 1085 2356 1090
rect 2406 1085 2754 1138
rect 3482 1098 3828 1138
rect 2350 1043 2754 1085
rect 3428 1046 3434 1098
rect 3486 1046 3828 1098
rect 2350 1038 2356 1043
rect 2406 1006 2754 1043
rect 2406 966 2466 1006
rect 2654 966 2754 1006
rect 3482 1024 3828 1046
rect 3482 972 3538 1024
rect 3732 972 3828 1024
rect 3482 966 3828 972
rect 2406 950 2754 966
rect 2192 850 2586 898
rect 3241 854 3693 914
rect 2192 276 2248 850
rect 2292 731 2298 783
rect 2350 778 2356 783
rect 2350 736 2526 778
rect 2350 731 2356 736
rect 2584 506 2824 538
rect 2192 228 2596 276
rect 2192 128 2248 228
rect 2792 164 2824 506
rect 3241 278 3301 854
rect 3334 706 3340 758
rect 3392 756 3398 758
rect 3436 756 3618 760
rect 3392 712 3618 756
rect 3392 708 3486 712
rect 3392 706 3398 708
rect 3669 472 3957 514
rect 3241 218 3685 278
rect 3241 182 3301 218
rect 3217 176 3301 182
rect 2957 164 3301 176
rect 326 79 468 82
rect -309 36 -303 41
rect 541 -20 671 40
rect 375 -46 671 -20
rect -571 -146 -103 -94
rect -567 -412 -515 -146
rect 375 -218 617 -46
rect 659 -218 671 -46
rect 375 -220 671 -218
rect -367 -310 -361 -258
rect -309 -263 -303 -258
rect -309 -305 -180 -263
rect -309 -310 -303 -305
rect -123 -306 71 -262
rect -567 -464 -115 -412
rect 25 -514 69 -306
rect 541 -314 671 -220
rect 729 -399 767 -105
rect 884 -108 922 82
rect 1651 80 2248 128
rect 2790 126 3301 164
rect 2790 116 3060 126
rect 1296 40 1694 80
rect 1939 78 1975 80
rect 1044 -164 1082 -120
rect 894 -280 934 -168
rect 1037 -170 1089 -164
rect 992 -194 996 -188
rect 1037 -228 1089 -222
rect 1296 -212 1336 40
rect 2192 -48 2248 80
rect 2384 44 2390 96
rect 2442 86 2448 96
rect 2792 86 2824 116
rect 2442 54 2824 86
rect 2957 80 3060 116
rect 2442 44 2448 54
rect 2192 -96 2598 -48
rect 2196 -104 2598 -96
rect 1296 -230 1338 -212
rect 1298 -280 1338 -230
rect 894 -320 1338 -280
rect 2198 -368 2256 -104
rect 2384 -248 2390 -196
rect 2442 -206 2448 -196
rect 2442 -238 2534 -206
rect 2442 -248 2448 -238
rect 2590 -256 2762 -216
rect 1037 -392 1089 -386
rect 729 -437 1037 -399
rect -329 -526 69 -514
rect -329 -566 -233 -526
rect -63 -566 69 -526
rect 888 -562 932 -437
rect 2198 -424 2602 -368
rect 1037 -450 1089 -444
rect 2710 -474 2750 -256
rect 2396 -490 2750 -474
rect 2396 -526 2476 -490
rect 2650 -514 2750 -490
rect 2650 -526 2748 -514
rect -329 -578 69 -566
rect -329 -630 27 -578
rect 2396 -606 2748 -526
rect -253 -828 -53 -630
rect 2462 -754 2662 -606
rect 3010 -939 3060 80
rect 3241 -124 3301 126
rect 3914 134 3956 472
rect 4041 134 4093 2586
rect 6495 2433 6553 2857
rect 6980 2706 7700 2750
rect 6980 2504 7024 2706
rect 7260 2580 7420 2664
rect 7130 2549 7188 2572
rect 6808 2210 6848 2446
rect 7130 2436 7188 2491
rect 7260 2380 7592 2580
rect 7656 2541 7700 2706
rect 7656 2487 8010 2541
rect 7260 2324 7420 2380
rect 5777 2170 6848 2210
rect 7656 2200 7700 2487
rect 4800 926 4862 1054
rect 4520 866 5144 926
rect 5204 866 5210 926
rect 4520 494 4580 866
rect 5060 764 5614 800
rect 5060 558 5096 764
rect 5258 646 5430 702
rect 5258 642 5546 646
rect 5144 606 5204 612
rect 5144 500 5204 546
rect 4790 243 4826 500
rect 5258 420 5268 642
rect 5314 446 5546 642
rect 5314 420 5430 446
rect 5258 360 5430 420
rect 5578 326 5614 764
rect 5777 326 5817 2170
rect 6522 2006 6604 2074
rect 6336 1994 6604 2006
rect 6336 1818 6550 1994
rect 6590 1818 6604 1994
rect 6336 1806 6604 1818
rect 6522 1722 6604 1806
rect 6652 1664 6693 1936
rect 6808 1920 6848 2170
rect 7178 2156 7700 2200
rect 6816 1774 6860 1872
rect 6956 1870 7012 1930
rect 6956 1808 7012 1814
rect 7178 1774 7222 2156
rect 6816 1730 7222 1774
rect 6644 1608 6956 1664
rect 7012 1608 7018 1664
rect 6780 1480 6850 1608
rect 6009 1115 6015 1167
rect 6067 1160 6073 1167
rect 6202 1166 6402 1478
rect 6130 1160 6494 1166
rect 6067 1122 6494 1160
rect 7216 1156 7416 1434
rect 7144 1154 7512 1156
rect 6067 1115 6073 1122
rect 6130 1102 6494 1122
rect 6984 1102 6990 1154
rect 7042 1102 7512 1154
rect 6130 1034 6228 1102
rect 6410 1034 6494 1102
rect 6130 1028 6494 1034
rect 7144 1054 7512 1102
rect 7144 994 7229 1054
rect 7423 994 7512 1054
rect 7144 984 7512 994
rect 5933 918 6349 974
rect 5933 784 5989 918
rect 6860 896 7364 956
rect 5933 658 5981 784
rect 6015 744 6067 750
rect 6067 699 6294 737
rect 6015 686 6067 692
rect 6860 668 6920 896
rect 6984 712 6990 764
rect 7042 712 7296 764
rect 5933 342 5989 658
rect 6350 596 6602 646
rect 6860 608 7066 668
rect 5933 326 6363 342
rect 5576 290 6363 326
rect 5222 286 6363 290
rect 5222 280 6003 286
rect 5222 254 5614 280
rect 3914 82 4093 134
rect 4262 193 4832 243
rect 3477 10 3483 62
rect 3535 57 3541 62
rect 3914 57 3956 82
rect 3535 15 3956 57
rect 3535 10 3541 15
rect 3241 -184 3705 -124
rect 3241 -446 3301 -184
rect 3477 -326 3483 -274
rect 3535 -279 3541 -274
rect 3535 -321 3638 -279
rect 3535 -326 3541 -321
rect 3684 -336 3862 -288
rect 3241 -506 3703 -446
rect 3814 -554 3862 -336
rect 3467 -560 3862 -554
rect 3467 -610 3549 -560
rect 3767 -610 3862 -560
rect 3467 -620 3862 -610
rect 3467 -674 3845 -620
rect 3589 -838 3789 -674
rect 4262 -939 4312 193
rect 4516 86 4634 158
rect 4516 68 4582 86
rect 4368 -108 4582 68
rect 4624 -108 4634 86
rect 4368 -132 4634 -108
rect 4516 -202 4634 -132
rect 4686 -260 4736 12
rect 4790 8 4826 193
rect 5002 -52 5050 8
rect 4846 -170 4882 -52
rect 5000 -58 5052 -52
rect 5000 -116 5052 -110
rect 5002 -122 5050 -116
rect 5222 -170 5258 254
rect 4846 -206 5258 -170
rect 5933 10 5989 280
rect 6551 270 6601 596
rect 7006 306 7066 608
rect 7354 536 7644 588
rect 7004 284 7368 306
rect 6856 270 7368 284
rect 6551 246 7368 270
rect 6551 230 7066 246
rect 6551 224 6906 230
rect 6090 122 6096 174
rect 6148 173 6154 174
rect 6551 173 6601 224
rect 6148 123 6601 173
rect 6148 122 6154 123
rect 5933 -46 6359 10
rect 4684 -312 4736 -260
rect 4994 -298 5000 -246
rect 5052 -298 5058 -246
rect 4684 -342 4732 -312
rect 5002 -342 5050 -298
rect 4684 -390 5050 -342
rect 5933 -322 5989 -46
rect 6096 -164 6148 -158
rect 6148 -215 6295 -165
rect 6096 -222 6148 -216
rect 6338 -228 6560 -172
rect 5933 -378 6351 -322
rect 4710 -458 5020 -390
rect 6504 -416 6560 -228
rect 6136 -428 6560 -416
rect 4772 -634 4972 -458
rect 6136 -476 6241 -428
rect 6407 -476 6560 -428
rect 6136 -508 6560 -476
rect 6136 -572 6504 -508
rect 6272 -732 6472 -572
rect 3010 -989 4312 -939
rect 6753 -904 6797 224
rect 7004 -54 7064 230
rect 7592 222 7644 536
rect 7956 222 8010 2487
rect 8096 222 8150 3811
rect 7592 168 8484 222
rect 7592 126 7644 168
rect 7118 74 7124 126
rect 7176 74 7644 126
rect 7839 -50 8321 -6
rect 6990 -114 7356 -54
rect 7004 -378 7064 -114
rect 7118 -274 7124 -222
rect 7176 -274 7306 -222
rect 7358 -330 7530 -292
rect 7004 -380 7220 -378
rect 7004 -428 7370 -380
rect 7492 -490 7530 -330
rect 7138 -500 7530 -490
rect 7138 -544 7241 -500
rect 7413 -544 7530 -500
rect 7138 -549 7530 -544
rect 7138 -616 7518 -549
rect 7238 -852 7438 -616
rect 7839 -904 7883 -50
rect 6753 -948 7883 -904
<< via1 >>
rect 3069 2964 3121 3016
rect 3069 2664 3121 2716
rect -447 1090 -395 1142
rect -447 781 -395 833
rect 7130 2857 7188 2915
rect 1056 536 1108 588
rect 1326 654 1378 706
rect -361 36 -309 88
rect 2916 1992 2968 2044
rect 2916 1748 2968 1800
rect 2298 1038 2350 1090
rect 3434 1046 3486 1098
rect 2298 731 2350 783
rect 3340 706 3392 758
rect -361 -310 -309 -258
rect 1037 -222 1089 -170
rect 2390 44 2442 96
rect 2390 -248 2442 -196
rect 1037 -444 1089 -392
rect 7130 2491 7188 2549
rect 5144 866 5204 926
rect 5144 546 5204 606
rect 6956 1814 7012 1870
rect 6956 1608 7012 1664
rect 6015 1115 6067 1167
rect 6990 1102 7042 1154
rect 6015 692 6067 744
rect 6990 712 7042 764
rect 3483 10 3535 62
rect 3483 -326 3535 -274
rect 5000 -110 5052 -58
rect 6096 122 6148 174
rect 5000 -298 5052 -246
rect 6096 -216 6148 -164
rect 7124 74 7176 126
rect 7124 -274 7176 -222
<< metal2 >>
rect 3063 2964 3069 3016
rect 3121 2964 3127 3016
rect 3075 2716 3115 2964
rect 7130 2915 7188 2921
rect 3063 2664 3069 2716
rect 3121 2664 3127 2716
rect 7130 2549 7188 2857
rect 7124 2491 7130 2549
rect 7188 2491 7194 2549
rect 2910 1992 2916 2044
rect 2968 1992 2974 2044
rect 2916 1800 2968 1992
rect 6950 1814 6956 1870
rect 7012 1814 7018 1870
rect 2916 1742 2968 1748
rect 6956 1664 7012 1814
rect 6956 1602 7012 1608
rect 6015 1167 6067 1173
rect -447 1142 -395 1148
rect 6015 1109 6067 1115
rect 6990 1154 7042 1160
rect 3434 1098 3486 1104
rect -447 1084 -395 1090
rect 2298 1090 2350 1096
rect -444 839 -398 1084
rect 2298 1032 2350 1038
rect 3342 1048 3434 1096
rect -447 833 -395 839
rect 2303 789 2345 1032
rect -447 775 -395 781
rect 2298 783 2350 789
rect 3342 764 3390 1048
rect 3434 1040 3486 1046
rect 5144 926 5204 932
rect 2298 725 2350 731
rect 3340 758 3392 764
rect 1320 700 1326 706
rect 1062 660 1326 700
rect 1062 588 1102 660
rect 1320 654 1326 660
rect 1378 654 1384 706
rect 3340 700 3392 706
rect 5144 606 5204 866
rect 6022 744 6060 1109
rect 6990 764 7042 1102
rect 6009 692 6015 744
rect 6067 692 6073 744
rect 6990 706 7042 712
rect 1050 536 1056 588
rect 1108 536 1114 588
rect 5138 546 5144 606
rect 5204 546 5210 606
rect 6096 174 6148 180
rect 6096 116 6148 122
rect 7124 126 7176 132
rect 2390 96 2442 102
rect -361 88 -309 94
rect 2390 38 2442 44
rect 3483 62 3535 68
rect -361 30 -309 36
rect -356 -252 -314 30
rect 1031 -222 1037 -170
rect 1089 -222 1095 -170
rect 2400 -190 2432 38
rect 3483 4 3535 10
rect 2390 -196 2442 -190
rect -361 -258 -309 -252
rect -361 -316 -309 -310
rect 1044 -392 1082 -222
rect 2390 -254 2442 -248
rect 3488 -268 3530 4
rect 4994 -110 5000 -58
rect 5052 -110 5058 -58
rect 5002 -240 5050 -110
rect 6097 -164 6147 116
rect 6090 -216 6096 -164
rect 6148 -216 6154 -164
rect 7124 -222 7176 74
rect 5000 -246 5052 -240
rect 3483 -274 3535 -268
rect 7124 -280 7176 -274
rect 5000 -304 5052 -298
rect 3483 -332 3535 -326
rect 1031 -444 1037 -392
rect 1089 -444 1095 -392
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM1
timestamp 1713377695
transform 1 0 2557 0 1 565
box -211 -469 211 469
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1713377695
transform 1 0 7329 0 1 -246
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM3
timestamp 1713377695
transform 0 -1 6851 1 0 2471
box -211 -469 211 469
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1713377695
transform 0 -1 4868 1 0 -23
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 1713377695
transform 1 0 2563 0 1 -238
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM6
timestamp 1713377695
transform 0 -1 919 1 0 433
box -211 -469 211 469
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM7
timestamp 1713377695
transform 0 1 2781 -1 0 2615
box -211 -469 211 469
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1713377695
transform 0 -1 2788 1 0 2047
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM9
timestamp 1713377695
transform 0 1 4859 -1 0 529
box -211 -469 211 469
use sky130_fd_pr__nfet_01v8_648S5X  XM10
timestamp 1713377695
transform 0 -1 6826 1 0 1897
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM11
timestamp 1713377695
transform 0 -1 908 1 0 -139
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM12
timestamp 1713377695
transform 1 0 3647 0 1 563
box -211 -469 211 469
use sky130_fd_pr__nfet_01v8_648S5X  XM13
timestamp 1713377695
transform 1 0 6325 0 1 -186
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM14
timestamp 1713377695
transform 1 0 7323 0 1 591
box -211 -469 211 469
use sky130_fd_pr__nfet_01v8_648S5X  XM15
timestamp 1713377695
transform 1 0 3659 0 1 -314
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM16
timestamp 1713377695
transform 1 0 -144 0 1 605
box -211 -469 211 469
use sky130_fd_pr__pfet_01v8_XJ7KDL  XM17
timestamp 1713377695
transform 1 0 6319 0 1 637
box -211 -469 211 469
use sky130_fd_pr__nfet_01v8_648S5X  XM18
timestamp 1713377695
transform 1 0 -148 0 1 -280
box -211 -310 211 310
<< labels >>
flabel metal1 263 152 263 152 0 FreeSans 320 0 0 0 clk_b
flabel metal1 -253 -828 -53 -628 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 -253 1246 -53 1446 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 375 -220 575 -20 0 FreeSans 256 90 0 0 GND
port 2 nsew
flabel metal1 1371 340 1571 540 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 8433 192 8433 192 0 FreeSans 320 0 0 0 q_b
flabel metal1 3589 -838 3789 -638 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 2462 -754 2662 -554 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 6814 1516 6814 1516 0 FreeSans 320 0 0 0 clk_b
flabel metal1 6754 3006 6954 3206 0 FreeSans 256 180 0 0 clk
port 3 nsew
flabel metal1 6336 1806 6536 2006 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 7392 2380 7592 2580 0 FreeSans 256 90 0 0 VDD
port 1 nsew
flabel metal1 7238 -852 7438 -652 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 7216 1234 7416 1434 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 6272 -732 6472 -532 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 6202 1278 6402 1478 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 908 -530 908 -530 0 FreeSans 320 0 0 0 clk_b
flabel metal1 802 940 1002 1140 0 FreeSans 256 180 0 0 clk
port 3 nsew
flabel metal1 5346 446 5546 646 0 FreeSans 256 90 0 0 VDD
port 1 nsew
flabel metal1 4368 -132 4568 68 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 4772 -634 4972 -434 0 FreeSans 256 0 0 0 clk
port 3 nsew
flabel metal1 4832 1030 4832 1030 0 FreeSans 320 0 0 0 clk_b
flabel metal1 3542 1184 3742 1384 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 2462 1146 2662 1346 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 2658 1484 2858 1684 0 FreeSans 256 0 0 0 clk
port 3 nsew
flabel metal1 2760 3072 2760 3072 0 FreeSans 480 0 0 0 clk_b
flabel metal1 2244 1958 2444 2158 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 3276 2522 3476 2722 0 FreeSans 256 90 0 0 VDD
port 1 nsew
flabel metal1 -833 162 -633 362 0 FreeSans 256 180 0 0 clk
port 3 nsew
<< end >>
