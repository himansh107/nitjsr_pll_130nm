magic
tech sky130A
magscale 1 2
timestamp 1714629389
<< metal3 >>
rect -39552 37772 -33180 37800
rect -39552 31748 -33264 37772
rect -33200 31748 -33180 37772
rect -39552 31720 -33180 31748
rect -32940 37772 -26568 37800
rect -32940 31748 -26652 37772
rect -26588 31748 -26568 37772
rect -32940 31720 -26568 31748
rect -26328 37772 -19956 37800
rect -26328 31748 -20040 37772
rect -19976 31748 -19956 37772
rect -26328 31720 -19956 31748
rect -19716 37772 -13344 37800
rect -19716 31748 -13428 37772
rect -13364 31748 -13344 37772
rect -19716 31720 -13344 31748
rect -13104 37772 -6732 37800
rect -13104 31748 -6816 37772
rect -6752 31748 -6732 37772
rect -13104 31720 -6732 31748
rect -6492 37772 -120 37800
rect -6492 31748 -204 37772
rect -140 31748 -120 37772
rect -6492 31720 -120 31748
rect 120 37772 6492 37800
rect 120 31748 6408 37772
rect 6472 31748 6492 37772
rect 120 31720 6492 31748
rect 6732 37772 13104 37800
rect 6732 31748 13020 37772
rect 13084 31748 13104 37772
rect 6732 31720 13104 31748
rect 13344 37772 19716 37800
rect 13344 31748 19632 37772
rect 19696 31748 19716 37772
rect 13344 31720 19716 31748
rect 19956 37772 26328 37800
rect 19956 31748 26244 37772
rect 26308 31748 26328 37772
rect 19956 31720 26328 31748
rect 26568 37772 32940 37800
rect 26568 31748 32856 37772
rect 32920 31748 32940 37772
rect 26568 31720 32940 31748
rect 33180 37772 39552 37800
rect 33180 31748 39468 37772
rect 39532 31748 39552 37772
rect 33180 31720 39552 31748
rect -39552 31452 -33180 31480
rect -39552 25428 -33264 31452
rect -33200 25428 -33180 31452
rect -39552 25400 -33180 25428
rect -32940 31452 -26568 31480
rect -32940 25428 -26652 31452
rect -26588 25428 -26568 31452
rect -32940 25400 -26568 25428
rect -26328 31452 -19956 31480
rect -26328 25428 -20040 31452
rect -19976 25428 -19956 31452
rect -26328 25400 -19956 25428
rect -19716 31452 -13344 31480
rect -19716 25428 -13428 31452
rect -13364 25428 -13344 31452
rect -19716 25400 -13344 25428
rect -13104 31452 -6732 31480
rect -13104 25428 -6816 31452
rect -6752 25428 -6732 31452
rect -13104 25400 -6732 25428
rect -6492 31452 -120 31480
rect -6492 25428 -204 31452
rect -140 25428 -120 31452
rect -6492 25400 -120 25428
rect 120 31452 6492 31480
rect 120 25428 6408 31452
rect 6472 25428 6492 31452
rect 120 25400 6492 25428
rect 6732 31452 13104 31480
rect 6732 25428 13020 31452
rect 13084 25428 13104 31452
rect 6732 25400 13104 25428
rect 13344 31452 19716 31480
rect 13344 25428 19632 31452
rect 19696 25428 19716 31452
rect 13344 25400 19716 25428
rect 19956 31452 26328 31480
rect 19956 25428 26244 31452
rect 26308 25428 26328 31452
rect 19956 25400 26328 25428
rect 26568 31452 32940 31480
rect 26568 25428 32856 31452
rect 32920 25428 32940 31452
rect 26568 25400 32940 25428
rect 33180 31452 39552 31480
rect 33180 25428 39468 31452
rect 39532 25428 39552 31452
rect 33180 25400 39552 25428
rect -39552 25132 -33180 25160
rect -39552 19108 -33264 25132
rect -33200 19108 -33180 25132
rect -39552 19080 -33180 19108
rect -32940 25132 -26568 25160
rect -32940 19108 -26652 25132
rect -26588 19108 -26568 25132
rect -32940 19080 -26568 19108
rect -26328 25132 -19956 25160
rect -26328 19108 -20040 25132
rect -19976 19108 -19956 25132
rect -26328 19080 -19956 19108
rect -19716 25132 -13344 25160
rect -19716 19108 -13428 25132
rect -13364 19108 -13344 25132
rect -19716 19080 -13344 19108
rect -13104 25132 -6732 25160
rect -13104 19108 -6816 25132
rect -6752 19108 -6732 25132
rect -13104 19080 -6732 19108
rect -6492 25132 -120 25160
rect -6492 19108 -204 25132
rect -140 19108 -120 25132
rect -6492 19080 -120 19108
rect 120 25132 6492 25160
rect 120 19108 6408 25132
rect 6472 19108 6492 25132
rect 120 19080 6492 19108
rect 6732 25132 13104 25160
rect 6732 19108 13020 25132
rect 13084 19108 13104 25132
rect 6732 19080 13104 19108
rect 13344 25132 19716 25160
rect 13344 19108 19632 25132
rect 19696 19108 19716 25132
rect 13344 19080 19716 19108
rect 19956 25132 26328 25160
rect 19956 19108 26244 25132
rect 26308 19108 26328 25132
rect 19956 19080 26328 19108
rect 26568 25132 32940 25160
rect 26568 19108 32856 25132
rect 32920 19108 32940 25132
rect 26568 19080 32940 19108
rect 33180 25132 39552 25160
rect 33180 19108 39468 25132
rect 39532 19108 39552 25132
rect 33180 19080 39552 19108
rect -39552 18812 -33180 18840
rect -39552 12788 -33264 18812
rect -33200 12788 -33180 18812
rect -39552 12760 -33180 12788
rect -32940 18812 -26568 18840
rect -32940 12788 -26652 18812
rect -26588 12788 -26568 18812
rect -32940 12760 -26568 12788
rect -26328 18812 -19956 18840
rect -26328 12788 -20040 18812
rect -19976 12788 -19956 18812
rect -26328 12760 -19956 12788
rect -19716 18812 -13344 18840
rect -19716 12788 -13428 18812
rect -13364 12788 -13344 18812
rect -19716 12760 -13344 12788
rect -13104 18812 -6732 18840
rect -13104 12788 -6816 18812
rect -6752 12788 -6732 18812
rect -13104 12760 -6732 12788
rect -6492 18812 -120 18840
rect -6492 12788 -204 18812
rect -140 12788 -120 18812
rect -6492 12760 -120 12788
rect 120 18812 6492 18840
rect 120 12788 6408 18812
rect 6472 12788 6492 18812
rect 120 12760 6492 12788
rect 6732 18812 13104 18840
rect 6732 12788 13020 18812
rect 13084 12788 13104 18812
rect 6732 12760 13104 12788
rect 13344 18812 19716 18840
rect 13344 12788 19632 18812
rect 19696 12788 19716 18812
rect 13344 12760 19716 12788
rect 19956 18812 26328 18840
rect 19956 12788 26244 18812
rect 26308 12788 26328 18812
rect 19956 12760 26328 12788
rect 26568 18812 32940 18840
rect 26568 12788 32856 18812
rect 32920 12788 32940 18812
rect 26568 12760 32940 12788
rect 33180 18812 39552 18840
rect 33180 12788 39468 18812
rect 39532 12788 39552 18812
rect 33180 12760 39552 12788
rect -39552 12492 -33180 12520
rect -39552 6468 -33264 12492
rect -33200 6468 -33180 12492
rect -39552 6440 -33180 6468
rect -32940 12492 -26568 12520
rect -32940 6468 -26652 12492
rect -26588 6468 -26568 12492
rect -32940 6440 -26568 6468
rect -26328 12492 -19956 12520
rect -26328 6468 -20040 12492
rect -19976 6468 -19956 12492
rect -26328 6440 -19956 6468
rect -19716 12492 -13344 12520
rect -19716 6468 -13428 12492
rect -13364 6468 -13344 12492
rect -19716 6440 -13344 6468
rect -13104 12492 -6732 12520
rect -13104 6468 -6816 12492
rect -6752 6468 -6732 12492
rect -13104 6440 -6732 6468
rect -6492 12492 -120 12520
rect -6492 6468 -204 12492
rect -140 6468 -120 12492
rect -6492 6440 -120 6468
rect 120 12492 6492 12520
rect 120 6468 6408 12492
rect 6472 6468 6492 12492
rect 120 6440 6492 6468
rect 6732 12492 13104 12520
rect 6732 6468 13020 12492
rect 13084 6468 13104 12492
rect 6732 6440 13104 6468
rect 13344 12492 19716 12520
rect 13344 6468 19632 12492
rect 19696 6468 19716 12492
rect 13344 6440 19716 6468
rect 19956 12492 26328 12520
rect 19956 6468 26244 12492
rect 26308 6468 26328 12492
rect 19956 6440 26328 6468
rect 26568 12492 32940 12520
rect 26568 6468 32856 12492
rect 32920 6468 32940 12492
rect 26568 6440 32940 6468
rect 33180 12492 39552 12520
rect 33180 6468 39468 12492
rect 39532 6468 39552 12492
rect 33180 6440 39552 6468
rect -39552 6172 -33180 6200
rect -39552 148 -33264 6172
rect -33200 148 -33180 6172
rect -39552 120 -33180 148
rect -32940 6172 -26568 6200
rect -32940 148 -26652 6172
rect -26588 148 -26568 6172
rect -32940 120 -26568 148
rect -26328 6172 -19956 6200
rect -26328 148 -20040 6172
rect -19976 148 -19956 6172
rect -26328 120 -19956 148
rect -19716 6172 -13344 6200
rect -19716 148 -13428 6172
rect -13364 148 -13344 6172
rect -19716 120 -13344 148
rect -13104 6172 -6732 6200
rect -13104 148 -6816 6172
rect -6752 148 -6732 6172
rect -13104 120 -6732 148
rect -6492 6172 -120 6200
rect -6492 148 -204 6172
rect -140 148 -120 6172
rect -6492 120 -120 148
rect 120 6172 6492 6200
rect 120 148 6408 6172
rect 6472 148 6492 6172
rect 120 120 6492 148
rect 6732 6172 13104 6200
rect 6732 148 13020 6172
rect 13084 148 13104 6172
rect 6732 120 13104 148
rect 13344 6172 19716 6200
rect 13344 148 19632 6172
rect 19696 148 19716 6172
rect 13344 120 19716 148
rect 19956 6172 26328 6200
rect 19956 148 26244 6172
rect 26308 148 26328 6172
rect 19956 120 26328 148
rect 26568 6172 32940 6200
rect 26568 148 32856 6172
rect 32920 148 32940 6172
rect 26568 120 32940 148
rect 33180 6172 39552 6200
rect 33180 148 39468 6172
rect 39532 148 39552 6172
rect 33180 120 39552 148
rect -39552 -148 -33180 -120
rect -39552 -6172 -33264 -148
rect -33200 -6172 -33180 -148
rect -39552 -6200 -33180 -6172
rect -32940 -148 -26568 -120
rect -32940 -6172 -26652 -148
rect -26588 -6172 -26568 -148
rect -32940 -6200 -26568 -6172
rect -26328 -148 -19956 -120
rect -26328 -6172 -20040 -148
rect -19976 -6172 -19956 -148
rect -26328 -6200 -19956 -6172
rect -19716 -148 -13344 -120
rect -19716 -6172 -13428 -148
rect -13364 -6172 -13344 -148
rect -19716 -6200 -13344 -6172
rect -13104 -148 -6732 -120
rect -13104 -6172 -6816 -148
rect -6752 -6172 -6732 -148
rect -13104 -6200 -6732 -6172
rect -6492 -148 -120 -120
rect -6492 -6172 -204 -148
rect -140 -6172 -120 -148
rect -6492 -6200 -120 -6172
rect 120 -148 6492 -120
rect 120 -6172 6408 -148
rect 6472 -6172 6492 -148
rect 120 -6200 6492 -6172
rect 6732 -148 13104 -120
rect 6732 -6172 13020 -148
rect 13084 -6172 13104 -148
rect 6732 -6200 13104 -6172
rect 13344 -148 19716 -120
rect 13344 -6172 19632 -148
rect 19696 -6172 19716 -148
rect 13344 -6200 19716 -6172
rect 19956 -148 26328 -120
rect 19956 -6172 26244 -148
rect 26308 -6172 26328 -148
rect 19956 -6200 26328 -6172
rect 26568 -148 32940 -120
rect 26568 -6172 32856 -148
rect 32920 -6172 32940 -148
rect 26568 -6200 32940 -6172
rect 33180 -148 39552 -120
rect 33180 -6172 39468 -148
rect 39532 -6172 39552 -148
rect 33180 -6200 39552 -6172
rect -39552 -6468 -33180 -6440
rect -39552 -12492 -33264 -6468
rect -33200 -12492 -33180 -6468
rect -39552 -12520 -33180 -12492
rect -32940 -6468 -26568 -6440
rect -32940 -12492 -26652 -6468
rect -26588 -12492 -26568 -6468
rect -32940 -12520 -26568 -12492
rect -26328 -6468 -19956 -6440
rect -26328 -12492 -20040 -6468
rect -19976 -12492 -19956 -6468
rect -26328 -12520 -19956 -12492
rect -19716 -6468 -13344 -6440
rect -19716 -12492 -13428 -6468
rect -13364 -12492 -13344 -6468
rect -19716 -12520 -13344 -12492
rect -13104 -6468 -6732 -6440
rect -13104 -12492 -6816 -6468
rect -6752 -12492 -6732 -6468
rect -13104 -12520 -6732 -12492
rect -6492 -6468 -120 -6440
rect -6492 -12492 -204 -6468
rect -140 -12492 -120 -6468
rect -6492 -12520 -120 -12492
rect 120 -6468 6492 -6440
rect 120 -12492 6408 -6468
rect 6472 -12492 6492 -6468
rect 120 -12520 6492 -12492
rect 6732 -6468 13104 -6440
rect 6732 -12492 13020 -6468
rect 13084 -12492 13104 -6468
rect 6732 -12520 13104 -12492
rect 13344 -6468 19716 -6440
rect 13344 -12492 19632 -6468
rect 19696 -12492 19716 -6468
rect 13344 -12520 19716 -12492
rect 19956 -6468 26328 -6440
rect 19956 -12492 26244 -6468
rect 26308 -12492 26328 -6468
rect 19956 -12520 26328 -12492
rect 26568 -6468 32940 -6440
rect 26568 -12492 32856 -6468
rect 32920 -12492 32940 -6468
rect 26568 -12520 32940 -12492
rect 33180 -6468 39552 -6440
rect 33180 -12492 39468 -6468
rect 39532 -12492 39552 -6468
rect 33180 -12520 39552 -12492
rect -39552 -12788 -33180 -12760
rect -39552 -18812 -33264 -12788
rect -33200 -18812 -33180 -12788
rect -39552 -18840 -33180 -18812
rect -32940 -12788 -26568 -12760
rect -32940 -18812 -26652 -12788
rect -26588 -18812 -26568 -12788
rect -32940 -18840 -26568 -18812
rect -26328 -12788 -19956 -12760
rect -26328 -18812 -20040 -12788
rect -19976 -18812 -19956 -12788
rect -26328 -18840 -19956 -18812
rect -19716 -12788 -13344 -12760
rect -19716 -18812 -13428 -12788
rect -13364 -18812 -13344 -12788
rect -19716 -18840 -13344 -18812
rect -13104 -12788 -6732 -12760
rect -13104 -18812 -6816 -12788
rect -6752 -18812 -6732 -12788
rect -13104 -18840 -6732 -18812
rect -6492 -12788 -120 -12760
rect -6492 -18812 -204 -12788
rect -140 -18812 -120 -12788
rect -6492 -18840 -120 -18812
rect 120 -12788 6492 -12760
rect 120 -18812 6408 -12788
rect 6472 -18812 6492 -12788
rect 120 -18840 6492 -18812
rect 6732 -12788 13104 -12760
rect 6732 -18812 13020 -12788
rect 13084 -18812 13104 -12788
rect 6732 -18840 13104 -18812
rect 13344 -12788 19716 -12760
rect 13344 -18812 19632 -12788
rect 19696 -18812 19716 -12788
rect 13344 -18840 19716 -18812
rect 19956 -12788 26328 -12760
rect 19956 -18812 26244 -12788
rect 26308 -18812 26328 -12788
rect 19956 -18840 26328 -18812
rect 26568 -12788 32940 -12760
rect 26568 -18812 32856 -12788
rect 32920 -18812 32940 -12788
rect 26568 -18840 32940 -18812
rect 33180 -12788 39552 -12760
rect 33180 -18812 39468 -12788
rect 39532 -18812 39552 -12788
rect 33180 -18840 39552 -18812
rect -39552 -19108 -33180 -19080
rect -39552 -25132 -33264 -19108
rect -33200 -25132 -33180 -19108
rect -39552 -25160 -33180 -25132
rect -32940 -19108 -26568 -19080
rect -32940 -25132 -26652 -19108
rect -26588 -25132 -26568 -19108
rect -32940 -25160 -26568 -25132
rect -26328 -19108 -19956 -19080
rect -26328 -25132 -20040 -19108
rect -19976 -25132 -19956 -19108
rect -26328 -25160 -19956 -25132
rect -19716 -19108 -13344 -19080
rect -19716 -25132 -13428 -19108
rect -13364 -25132 -13344 -19108
rect -19716 -25160 -13344 -25132
rect -13104 -19108 -6732 -19080
rect -13104 -25132 -6816 -19108
rect -6752 -25132 -6732 -19108
rect -13104 -25160 -6732 -25132
rect -6492 -19108 -120 -19080
rect -6492 -25132 -204 -19108
rect -140 -25132 -120 -19108
rect -6492 -25160 -120 -25132
rect 120 -19108 6492 -19080
rect 120 -25132 6408 -19108
rect 6472 -25132 6492 -19108
rect 120 -25160 6492 -25132
rect 6732 -19108 13104 -19080
rect 6732 -25132 13020 -19108
rect 13084 -25132 13104 -19108
rect 6732 -25160 13104 -25132
rect 13344 -19108 19716 -19080
rect 13344 -25132 19632 -19108
rect 19696 -25132 19716 -19108
rect 13344 -25160 19716 -25132
rect 19956 -19108 26328 -19080
rect 19956 -25132 26244 -19108
rect 26308 -25132 26328 -19108
rect 19956 -25160 26328 -25132
rect 26568 -19108 32940 -19080
rect 26568 -25132 32856 -19108
rect 32920 -25132 32940 -19108
rect 26568 -25160 32940 -25132
rect 33180 -19108 39552 -19080
rect 33180 -25132 39468 -19108
rect 39532 -25132 39552 -19108
rect 33180 -25160 39552 -25132
rect -39552 -25428 -33180 -25400
rect -39552 -31452 -33264 -25428
rect -33200 -31452 -33180 -25428
rect -39552 -31480 -33180 -31452
rect -32940 -25428 -26568 -25400
rect -32940 -31452 -26652 -25428
rect -26588 -31452 -26568 -25428
rect -32940 -31480 -26568 -31452
rect -26328 -25428 -19956 -25400
rect -26328 -31452 -20040 -25428
rect -19976 -31452 -19956 -25428
rect -26328 -31480 -19956 -31452
rect -19716 -25428 -13344 -25400
rect -19716 -31452 -13428 -25428
rect -13364 -31452 -13344 -25428
rect -19716 -31480 -13344 -31452
rect -13104 -25428 -6732 -25400
rect -13104 -31452 -6816 -25428
rect -6752 -31452 -6732 -25428
rect -13104 -31480 -6732 -31452
rect -6492 -25428 -120 -25400
rect -6492 -31452 -204 -25428
rect -140 -31452 -120 -25428
rect -6492 -31480 -120 -31452
rect 120 -25428 6492 -25400
rect 120 -31452 6408 -25428
rect 6472 -31452 6492 -25428
rect 120 -31480 6492 -31452
rect 6732 -25428 13104 -25400
rect 6732 -31452 13020 -25428
rect 13084 -31452 13104 -25428
rect 6732 -31480 13104 -31452
rect 13344 -25428 19716 -25400
rect 13344 -31452 19632 -25428
rect 19696 -31452 19716 -25428
rect 13344 -31480 19716 -31452
rect 19956 -25428 26328 -25400
rect 19956 -31452 26244 -25428
rect 26308 -31452 26328 -25428
rect 19956 -31480 26328 -31452
rect 26568 -25428 32940 -25400
rect 26568 -31452 32856 -25428
rect 32920 -31452 32940 -25428
rect 26568 -31480 32940 -31452
rect 33180 -25428 39552 -25400
rect 33180 -31452 39468 -25428
rect 39532 -31452 39552 -25428
rect 33180 -31480 39552 -31452
rect -39552 -31748 -33180 -31720
rect -39552 -37772 -33264 -31748
rect -33200 -37772 -33180 -31748
rect -39552 -37800 -33180 -37772
rect -32940 -31748 -26568 -31720
rect -32940 -37772 -26652 -31748
rect -26588 -37772 -26568 -31748
rect -32940 -37800 -26568 -37772
rect -26328 -31748 -19956 -31720
rect -26328 -37772 -20040 -31748
rect -19976 -37772 -19956 -31748
rect -26328 -37800 -19956 -37772
rect -19716 -31748 -13344 -31720
rect -19716 -37772 -13428 -31748
rect -13364 -37772 -13344 -31748
rect -19716 -37800 -13344 -37772
rect -13104 -31748 -6732 -31720
rect -13104 -37772 -6816 -31748
rect -6752 -37772 -6732 -31748
rect -13104 -37800 -6732 -37772
rect -6492 -31748 -120 -31720
rect -6492 -37772 -204 -31748
rect -140 -37772 -120 -31748
rect -6492 -37800 -120 -37772
rect 120 -31748 6492 -31720
rect 120 -37772 6408 -31748
rect 6472 -37772 6492 -31748
rect 120 -37800 6492 -37772
rect 6732 -31748 13104 -31720
rect 6732 -37772 13020 -31748
rect 13084 -37772 13104 -31748
rect 6732 -37800 13104 -37772
rect 13344 -31748 19716 -31720
rect 13344 -37772 19632 -31748
rect 19696 -37772 19716 -31748
rect 13344 -37800 19716 -37772
rect 19956 -31748 26328 -31720
rect 19956 -37772 26244 -31748
rect 26308 -37772 26328 -31748
rect 19956 -37800 26328 -37772
rect 26568 -31748 32940 -31720
rect 26568 -37772 32856 -31748
rect 32920 -37772 32940 -31748
rect 26568 -37800 32940 -37772
rect 33180 -31748 39552 -31720
rect 33180 -37772 39468 -31748
rect 39532 -37772 39552 -31748
rect 33180 -37800 39552 -37772
<< via3 >>
rect -33264 31748 -33200 37772
rect -26652 31748 -26588 37772
rect -20040 31748 -19976 37772
rect -13428 31748 -13364 37772
rect -6816 31748 -6752 37772
rect -204 31748 -140 37772
rect 6408 31748 6472 37772
rect 13020 31748 13084 37772
rect 19632 31748 19696 37772
rect 26244 31748 26308 37772
rect 32856 31748 32920 37772
rect 39468 31748 39532 37772
rect -33264 25428 -33200 31452
rect -26652 25428 -26588 31452
rect -20040 25428 -19976 31452
rect -13428 25428 -13364 31452
rect -6816 25428 -6752 31452
rect -204 25428 -140 31452
rect 6408 25428 6472 31452
rect 13020 25428 13084 31452
rect 19632 25428 19696 31452
rect 26244 25428 26308 31452
rect 32856 25428 32920 31452
rect 39468 25428 39532 31452
rect -33264 19108 -33200 25132
rect -26652 19108 -26588 25132
rect -20040 19108 -19976 25132
rect -13428 19108 -13364 25132
rect -6816 19108 -6752 25132
rect -204 19108 -140 25132
rect 6408 19108 6472 25132
rect 13020 19108 13084 25132
rect 19632 19108 19696 25132
rect 26244 19108 26308 25132
rect 32856 19108 32920 25132
rect 39468 19108 39532 25132
rect -33264 12788 -33200 18812
rect -26652 12788 -26588 18812
rect -20040 12788 -19976 18812
rect -13428 12788 -13364 18812
rect -6816 12788 -6752 18812
rect -204 12788 -140 18812
rect 6408 12788 6472 18812
rect 13020 12788 13084 18812
rect 19632 12788 19696 18812
rect 26244 12788 26308 18812
rect 32856 12788 32920 18812
rect 39468 12788 39532 18812
rect -33264 6468 -33200 12492
rect -26652 6468 -26588 12492
rect -20040 6468 -19976 12492
rect -13428 6468 -13364 12492
rect -6816 6468 -6752 12492
rect -204 6468 -140 12492
rect 6408 6468 6472 12492
rect 13020 6468 13084 12492
rect 19632 6468 19696 12492
rect 26244 6468 26308 12492
rect 32856 6468 32920 12492
rect 39468 6468 39532 12492
rect -33264 148 -33200 6172
rect -26652 148 -26588 6172
rect -20040 148 -19976 6172
rect -13428 148 -13364 6172
rect -6816 148 -6752 6172
rect -204 148 -140 6172
rect 6408 148 6472 6172
rect 13020 148 13084 6172
rect 19632 148 19696 6172
rect 26244 148 26308 6172
rect 32856 148 32920 6172
rect 39468 148 39532 6172
rect -33264 -6172 -33200 -148
rect -26652 -6172 -26588 -148
rect -20040 -6172 -19976 -148
rect -13428 -6172 -13364 -148
rect -6816 -6172 -6752 -148
rect -204 -6172 -140 -148
rect 6408 -6172 6472 -148
rect 13020 -6172 13084 -148
rect 19632 -6172 19696 -148
rect 26244 -6172 26308 -148
rect 32856 -6172 32920 -148
rect 39468 -6172 39532 -148
rect -33264 -12492 -33200 -6468
rect -26652 -12492 -26588 -6468
rect -20040 -12492 -19976 -6468
rect -13428 -12492 -13364 -6468
rect -6816 -12492 -6752 -6468
rect -204 -12492 -140 -6468
rect 6408 -12492 6472 -6468
rect 13020 -12492 13084 -6468
rect 19632 -12492 19696 -6468
rect 26244 -12492 26308 -6468
rect 32856 -12492 32920 -6468
rect 39468 -12492 39532 -6468
rect -33264 -18812 -33200 -12788
rect -26652 -18812 -26588 -12788
rect -20040 -18812 -19976 -12788
rect -13428 -18812 -13364 -12788
rect -6816 -18812 -6752 -12788
rect -204 -18812 -140 -12788
rect 6408 -18812 6472 -12788
rect 13020 -18812 13084 -12788
rect 19632 -18812 19696 -12788
rect 26244 -18812 26308 -12788
rect 32856 -18812 32920 -12788
rect 39468 -18812 39532 -12788
rect -33264 -25132 -33200 -19108
rect -26652 -25132 -26588 -19108
rect -20040 -25132 -19976 -19108
rect -13428 -25132 -13364 -19108
rect -6816 -25132 -6752 -19108
rect -204 -25132 -140 -19108
rect 6408 -25132 6472 -19108
rect 13020 -25132 13084 -19108
rect 19632 -25132 19696 -19108
rect 26244 -25132 26308 -19108
rect 32856 -25132 32920 -19108
rect 39468 -25132 39532 -19108
rect -33264 -31452 -33200 -25428
rect -26652 -31452 -26588 -25428
rect -20040 -31452 -19976 -25428
rect -13428 -31452 -13364 -25428
rect -6816 -31452 -6752 -25428
rect -204 -31452 -140 -25428
rect 6408 -31452 6472 -25428
rect 13020 -31452 13084 -25428
rect 19632 -31452 19696 -25428
rect 26244 -31452 26308 -25428
rect 32856 -31452 32920 -25428
rect 39468 -31452 39532 -25428
rect -33264 -37772 -33200 -31748
rect -26652 -37772 -26588 -31748
rect -20040 -37772 -19976 -31748
rect -13428 -37772 -13364 -31748
rect -6816 -37772 -6752 -31748
rect -204 -37772 -140 -31748
rect 6408 -37772 6472 -31748
rect 13020 -37772 13084 -31748
rect 19632 -37772 19696 -31748
rect 26244 -37772 26308 -31748
rect 32856 -37772 32920 -31748
rect 39468 -37772 39532 -31748
<< mimcap >>
rect -39512 37720 -33512 37760
rect -39512 31800 -39472 37720
rect -33552 31800 -33512 37720
rect -39512 31760 -33512 31800
rect -32900 37720 -26900 37760
rect -32900 31800 -32860 37720
rect -26940 31800 -26900 37720
rect -32900 31760 -26900 31800
rect -26288 37720 -20288 37760
rect -26288 31800 -26248 37720
rect -20328 31800 -20288 37720
rect -26288 31760 -20288 31800
rect -19676 37720 -13676 37760
rect -19676 31800 -19636 37720
rect -13716 31800 -13676 37720
rect -19676 31760 -13676 31800
rect -13064 37720 -7064 37760
rect -13064 31800 -13024 37720
rect -7104 31800 -7064 37720
rect -13064 31760 -7064 31800
rect -6452 37720 -452 37760
rect -6452 31800 -6412 37720
rect -492 31800 -452 37720
rect -6452 31760 -452 31800
rect 160 37720 6160 37760
rect 160 31800 200 37720
rect 6120 31800 6160 37720
rect 160 31760 6160 31800
rect 6772 37720 12772 37760
rect 6772 31800 6812 37720
rect 12732 31800 12772 37720
rect 6772 31760 12772 31800
rect 13384 37720 19384 37760
rect 13384 31800 13424 37720
rect 19344 31800 19384 37720
rect 13384 31760 19384 31800
rect 19996 37720 25996 37760
rect 19996 31800 20036 37720
rect 25956 31800 25996 37720
rect 19996 31760 25996 31800
rect 26608 37720 32608 37760
rect 26608 31800 26648 37720
rect 32568 31800 32608 37720
rect 26608 31760 32608 31800
rect 33220 37720 39220 37760
rect 33220 31800 33260 37720
rect 39180 31800 39220 37720
rect 33220 31760 39220 31800
rect -39512 31400 -33512 31440
rect -39512 25480 -39472 31400
rect -33552 25480 -33512 31400
rect -39512 25440 -33512 25480
rect -32900 31400 -26900 31440
rect -32900 25480 -32860 31400
rect -26940 25480 -26900 31400
rect -32900 25440 -26900 25480
rect -26288 31400 -20288 31440
rect -26288 25480 -26248 31400
rect -20328 25480 -20288 31400
rect -26288 25440 -20288 25480
rect -19676 31400 -13676 31440
rect -19676 25480 -19636 31400
rect -13716 25480 -13676 31400
rect -19676 25440 -13676 25480
rect -13064 31400 -7064 31440
rect -13064 25480 -13024 31400
rect -7104 25480 -7064 31400
rect -13064 25440 -7064 25480
rect -6452 31400 -452 31440
rect -6452 25480 -6412 31400
rect -492 25480 -452 31400
rect -6452 25440 -452 25480
rect 160 31400 6160 31440
rect 160 25480 200 31400
rect 6120 25480 6160 31400
rect 160 25440 6160 25480
rect 6772 31400 12772 31440
rect 6772 25480 6812 31400
rect 12732 25480 12772 31400
rect 6772 25440 12772 25480
rect 13384 31400 19384 31440
rect 13384 25480 13424 31400
rect 19344 25480 19384 31400
rect 13384 25440 19384 25480
rect 19996 31400 25996 31440
rect 19996 25480 20036 31400
rect 25956 25480 25996 31400
rect 19996 25440 25996 25480
rect 26608 31400 32608 31440
rect 26608 25480 26648 31400
rect 32568 25480 32608 31400
rect 26608 25440 32608 25480
rect 33220 31400 39220 31440
rect 33220 25480 33260 31400
rect 39180 25480 39220 31400
rect 33220 25440 39220 25480
rect -39512 25080 -33512 25120
rect -39512 19160 -39472 25080
rect -33552 19160 -33512 25080
rect -39512 19120 -33512 19160
rect -32900 25080 -26900 25120
rect -32900 19160 -32860 25080
rect -26940 19160 -26900 25080
rect -32900 19120 -26900 19160
rect -26288 25080 -20288 25120
rect -26288 19160 -26248 25080
rect -20328 19160 -20288 25080
rect -26288 19120 -20288 19160
rect -19676 25080 -13676 25120
rect -19676 19160 -19636 25080
rect -13716 19160 -13676 25080
rect -19676 19120 -13676 19160
rect -13064 25080 -7064 25120
rect -13064 19160 -13024 25080
rect -7104 19160 -7064 25080
rect -13064 19120 -7064 19160
rect -6452 25080 -452 25120
rect -6452 19160 -6412 25080
rect -492 19160 -452 25080
rect -6452 19120 -452 19160
rect 160 25080 6160 25120
rect 160 19160 200 25080
rect 6120 19160 6160 25080
rect 160 19120 6160 19160
rect 6772 25080 12772 25120
rect 6772 19160 6812 25080
rect 12732 19160 12772 25080
rect 6772 19120 12772 19160
rect 13384 25080 19384 25120
rect 13384 19160 13424 25080
rect 19344 19160 19384 25080
rect 13384 19120 19384 19160
rect 19996 25080 25996 25120
rect 19996 19160 20036 25080
rect 25956 19160 25996 25080
rect 19996 19120 25996 19160
rect 26608 25080 32608 25120
rect 26608 19160 26648 25080
rect 32568 19160 32608 25080
rect 26608 19120 32608 19160
rect 33220 25080 39220 25120
rect 33220 19160 33260 25080
rect 39180 19160 39220 25080
rect 33220 19120 39220 19160
rect -39512 18760 -33512 18800
rect -39512 12840 -39472 18760
rect -33552 12840 -33512 18760
rect -39512 12800 -33512 12840
rect -32900 18760 -26900 18800
rect -32900 12840 -32860 18760
rect -26940 12840 -26900 18760
rect -32900 12800 -26900 12840
rect -26288 18760 -20288 18800
rect -26288 12840 -26248 18760
rect -20328 12840 -20288 18760
rect -26288 12800 -20288 12840
rect -19676 18760 -13676 18800
rect -19676 12840 -19636 18760
rect -13716 12840 -13676 18760
rect -19676 12800 -13676 12840
rect -13064 18760 -7064 18800
rect -13064 12840 -13024 18760
rect -7104 12840 -7064 18760
rect -13064 12800 -7064 12840
rect -6452 18760 -452 18800
rect -6452 12840 -6412 18760
rect -492 12840 -452 18760
rect -6452 12800 -452 12840
rect 160 18760 6160 18800
rect 160 12840 200 18760
rect 6120 12840 6160 18760
rect 160 12800 6160 12840
rect 6772 18760 12772 18800
rect 6772 12840 6812 18760
rect 12732 12840 12772 18760
rect 6772 12800 12772 12840
rect 13384 18760 19384 18800
rect 13384 12840 13424 18760
rect 19344 12840 19384 18760
rect 13384 12800 19384 12840
rect 19996 18760 25996 18800
rect 19996 12840 20036 18760
rect 25956 12840 25996 18760
rect 19996 12800 25996 12840
rect 26608 18760 32608 18800
rect 26608 12840 26648 18760
rect 32568 12840 32608 18760
rect 26608 12800 32608 12840
rect 33220 18760 39220 18800
rect 33220 12840 33260 18760
rect 39180 12840 39220 18760
rect 33220 12800 39220 12840
rect -39512 12440 -33512 12480
rect -39512 6520 -39472 12440
rect -33552 6520 -33512 12440
rect -39512 6480 -33512 6520
rect -32900 12440 -26900 12480
rect -32900 6520 -32860 12440
rect -26940 6520 -26900 12440
rect -32900 6480 -26900 6520
rect -26288 12440 -20288 12480
rect -26288 6520 -26248 12440
rect -20328 6520 -20288 12440
rect -26288 6480 -20288 6520
rect -19676 12440 -13676 12480
rect -19676 6520 -19636 12440
rect -13716 6520 -13676 12440
rect -19676 6480 -13676 6520
rect -13064 12440 -7064 12480
rect -13064 6520 -13024 12440
rect -7104 6520 -7064 12440
rect -13064 6480 -7064 6520
rect -6452 12440 -452 12480
rect -6452 6520 -6412 12440
rect -492 6520 -452 12440
rect -6452 6480 -452 6520
rect 160 12440 6160 12480
rect 160 6520 200 12440
rect 6120 6520 6160 12440
rect 160 6480 6160 6520
rect 6772 12440 12772 12480
rect 6772 6520 6812 12440
rect 12732 6520 12772 12440
rect 6772 6480 12772 6520
rect 13384 12440 19384 12480
rect 13384 6520 13424 12440
rect 19344 6520 19384 12440
rect 13384 6480 19384 6520
rect 19996 12440 25996 12480
rect 19996 6520 20036 12440
rect 25956 6520 25996 12440
rect 19996 6480 25996 6520
rect 26608 12440 32608 12480
rect 26608 6520 26648 12440
rect 32568 6520 32608 12440
rect 26608 6480 32608 6520
rect 33220 12440 39220 12480
rect 33220 6520 33260 12440
rect 39180 6520 39220 12440
rect 33220 6480 39220 6520
rect -39512 6120 -33512 6160
rect -39512 200 -39472 6120
rect -33552 200 -33512 6120
rect -39512 160 -33512 200
rect -32900 6120 -26900 6160
rect -32900 200 -32860 6120
rect -26940 200 -26900 6120
rect -32900 160 -26900 200
rect -26288 6120 -20288 6160
rect -26288 200 -26248 6120
rect -20328 200 -20288 6120
rect -26288 160 -20288 200
rect -19676 6120 -13676 6160
rect -19676 200 -19636 6120
rect -13716 200 -13676 6120
rect -19676 160 -13676 200
rect -13064 6120 -7064 6160
rect -13064 200 -13024 6120
rect -7104 200 -7064 6120
rect -13064 160 -7064 200
rect -6452 6120 -452 6160
rect -6452 200 -6412 6120
rect -492 200 -452 6120
rect -6452 160 -452 200
rect 160 6120 6160 6160
rect 160 200 200 6120
rect 6120 200 6160 6120
rect 160 160 6160 200
rect 6772 6120 12772 6160
rect 6772 200 6812 6120
rect 12732 200 12772 6120
rect 6772 160 12772 200
rect 13384 6120 19384 6160
rect 13384 200 13424 6120
rect 19344 200 19384 6120
rect 13384 160 19384 200
rect 19996 6120 25996 6160
rect 19996 200 20036 6120
rect 25956 200 25996 6120
rect 19996 160 25996 200
rect 26608 6120 32608 6160
rect 26608 200 26648 6120
rect 32568 200 32608 6120
rect 26608 160 32608 200
rect 33220 6120 39220 6160
rect 33220 200 33260 6120
rect 39180 200 39220 6120
rect 33220 160 39220 200
rect -39512 -200 -33512 -160
rect -39512 -6120 -39472 -200
rect -33552 -6120 -33512 -200
rect -39512 -6160 -33512 -6120
rect -32900 -200 -26900 -160
rect -32900 -6120 -32860 -200
rect -26940 -6120 -26900 -200
rect -32900 -6160 -26900 -6120
rect -26288 -200 -20288 -160
rect -26288 -6120 -26248 -200
rect -20328 -6120 -20288 -200
rect -26288 -6160 -20288 -6120
rect -19676 -200 -13676 -160
rect -19676 -6120 -19636 -200
rect -13716 -6120 -13676 -200
rect -19676 -6160 -13676 -6120
rect -13064 -200 -7064 -160
rect -13064 -6120 -13024 -200
rect -7104 -6120 -7064 -200
rect -13064 -6160 -7064 -6120
rect -6452 -200 -452 -160
rect -6452 -6120 -6412 -200
rect -492 -6120 -452 -200
rect -6452 -6160 -452 -6120
rect 160 -200 6160 -160
rect 160 -6120 200 -200
rect 6120 -6120 6160 -200
rect 160 -6160 6160 -6120
rect 6772 -200 12772 -160
rect 6772 -6120 6812 -200
rect 12732 -6120 12772 -200
rect 6772 -6160 12772 -6120
rect 13384 -200 19384 -160
rect 13384 -6120 13424 -200
rect 19344 -6120 19384 -200
rect 13384 -6160 19384 -6120
rect 19996 -200 25996 -160
rect 19996 -6120 20036 -200
rect 25956 -6120 25996 -200
rect 19996 -6160 25996 -6120
rect 26608 -200 32608 -160
rect 26608 -6120 26648 -200
rect 32568 -6120 32608 -200
rect 26608 -6160 32608 -6120
rect 33220 -200 39220 -160
rect 33220 -6120 33260 -200
rect 39180 -6120 39220 -200
rect 33220 -6160 39220 -6120
rect -39512 -6520 -33512 -6480
rect -39512 -12440 -39472 -6520
rect -33552 -12440 -33512 -6520
rect -39512 -12480 -33512 -12440
rect -32900 -6520 -26900 -6480
rect -32900 -12440 -32860 -6520
rect -26940 -12440 -26900 -6520
rect -32900 -12480 -26900 -12440
rect -26288 -6520 -20288 -6480
rect -26288 -12440 -26248 -6520
rect -20328 -12440 -20288 -6520
rect -26288 -12480 -20288 -12440
rect -19676 -6520 -13676 -6480
rect -19676 -12440 -19636 -6520
rect -13716 -12440 -13676 -6520
rect -19676 -12480 -13676 -12440
rect -13064 -6520 -7064 -6480
rect -13064 -12440 -13024 -6520
rect -7104 -12440 -7064 -6520
rect -13064 -12480 -7064 -12440
rect -6452 -6520 -452 -6480
rect -6452 -12440 -6412 -6520
rect -492 -12440 -452 -6520
rect -6452 -12480 -452 -12440
rect 160 -6520 6160 -6480
rect 160 -12440 200 -6520
rect 6120 -12440 6160 -6520
rect 160 -12480 6160 -12440
rect 6772 -6520 12772 -6480
rect 6772 -12440 6812 -6520
rect 12732 -12440 12772 -6520
rect 6772 -12480 12772 -12440
rect 13384 -6520 19384 -6480
rect 13384 -12440 13424 -6520
rect 19344 -12440 19384 -6520
rect 13384 -12480 19384 -12440
rect 19996 -6520 25996 -6480
rect 19996 -12440 20036 -6520
rect 25956 -12440 25996 -6520
rect 19996 -12480 25996 -12440
rect 26608 -6520 32608 -6480
rect 26608 -12440 26648 -6520
rect 32568 -12440 32608 -6520
rect 26608 -12480 32608 -12440
rect 33220 -6520 39220 -6480
rect 33220 -12440 33260 -6520
rect 39180 -12440 39220 -6520
rect 33220 -12480 39220 -12440
rect -39512 -12840 -33512 -12800
rect -39512 -18760 -39472 -12840
rect -33552 -18760 -33512 -12840
rect -39512 -18800 -33512 -18760
rect -32900 -12840 -26900 -12800
rect -32900 -18760 -32860 -12840
rect -26940 -18760 -26900 -12840
rect -32900 -18800 -26900 -18760
rect -26288 -12840 -20288 -12800
rect -26288 -18760 -26248 -12840
rect -20328 -18760 -20288 -12840
rect -26288 -18800 -20288 -18760
rect -19676 -12840 -13676 -12800
rect -19676 -18760 -19636 -12840
rect -13716 -18760 -13676 -12840
rect -19676 -18800 -13676 -18760
rect -13064 -12840 -7064 -12800
rect -13064 -18760 -13024 -12840
rect -7104 -18760 -7064 -12840
rect -13064 -18800 -7064 -18760
rect -6452 -12840 -452 -12800
rect -6452 -18760 -6412 -12840
rect -492 -18760 -452 -12840
rect -6452 -18800 -452 -18760
rect 160 -12840 6160 -12800
rect 160 -18760 200 -12840
rect 6120 -18760 6160 -12840
rect 160 -18800 6160 -18760
rect 6772 -12840 12772 -12800
rect 6772 -18760 6812 -12840
rect 12732 -18760 12772 -12840
rect 6772 -18800 12772 -18760
rect 13384 -12840 19384 -12800
rect 13384 -18760 13424 -12840
rect 19344 -18760 19384 -12840
rect 13384 -18800 19384 -18760
rect 19996 -12840 25996 -12800
rect 19996 -18760 20036 -12840
rect 25956 -18760 25996 -12840
rect 19996 -18800 25996 -18760
rect 26608 -12840 32608 -12800
rect 26608 -18760 26648 -12840
rect 32568 -18760 32608 -12840
rect 26608 -18800 32608 -18760
rect 33220 -12840 39220 -12800
rect 33220 -18760 33260 -12840
rect 39180 -18760 39220 -12840
rect 33220 -18800 39220 -18760
rect -39512 -19160 -33512 -19120
rect -39512 -25080 -39472 -19160
rect -33552 -25080 -33512 -19160
rect -39512 -25120 -33512 -25080
rect -32900 -19160 -26900 -19120
rect -32900 -25080 -32860 -19160
rect -26940 -25080 -26900 -19160
rect -32900 -25120 -26900 -25080
rect -26288 -19160 -20288 -19120
rect -26288 -25080 -26248 -19160
rect -20328 -25080 -20288 -19160
rect -26288 -25120 -20288 -25080
rect -19676 -19160 -13676 -19120
rect -19676 -25080 -19636 -19160
rect -13716 -25080 -13676 -19160
rect -19676 -25120 -13676 -25080
rect -13064 -19160 -7064 -19120
rect -13064 -25080 -13024 -19160
rect -7104 -25080 -7064 -19160
rect -13064 -25120 -7064 -25080
rect -6452 -19160 -452 -19120
rect -6452 -25080 -6412 -19160
rect -492 -25080 -452 -19160
rect -6452 -25120 -452 -25080
rect 160 -19160 6160 -19120
rect 160 -25080 200 -19160
rect 6120 -25080 6160 -19160
rect 160 -25120 6160 -25080
rect 6772 -19160 12772 -19120
rect 6772 -25080 6812 -19160
rect 12732 -25080 12772 -19160
rect 6772 -25120 12772 -25080
rect 13384 -19160 19384 -19120
rect 13384 -25080 13424 -19160
rect 19344 -25080 19384 -19160
rect 13384 -25120 19384 -25080
rect 19996 -19160 25996 -19120
rect 19996 -25080 20036 -19160
rect 25956 -25080 25996 -19160
rect 19996 -25120 25996 -25080
rect 26608 -19160 32608 -19120
rect 26608 -25080 26648 -19160
rect 32568 -25080 32608 -19160
rect 26608 -25120 32608 -25080
rect 33220 -19160 39220 -19120
rect 33220 -25080 33260 -19160
rect 39180 -25080 39220 -19160
rect 33220 -25120 39220 -25080
rect -39512 -25480 -33512 -25440
rect -39512 -31400 -39472 -25480
rect -33552 -31400 -33512 -25480
rect -39512 -31440 -33512 -31400
rect -32900 -25480 -26900 -25440
rect -32900 -31400 -32860 -25480
rect -26940 -31400 -26900 -25480
rect -32900 -31440 -26900 -31400
rect -26288 -25480 -20288 -25440
rect -26288 -31400 -26248 -25480
rect -20328 -31400 -20288 -25480
rect -26288 -31440 -20288 -31400
rect -19676 -25480 -13676 -25440
rect -19676 -31400 -19636 -25480
rect -13716 -31400 -13676 -25480
rect -19676 -31440 -13676 -31400
rect -13064 -25480 -7064 -25440
rect -13064 -31400 -13024 -25480
rect -7104 -31400 -7064 -25480
rect -13064 -31440 -7064 -31400
rect -6452 -25480 -452 -25440
rect -6452 -31400 -6412 -25480
rect -492 -31400 -452 -25480
rect -6452 -31440 -452 -31400
rect 160 -25480 6160 -25440
rect 160 -31400 200 -25480
rect 6120 -31400 6160 -25480
rect 160 -31440 6160 -31400
rect 6772 -25480 12772 -25440
rect 6772 -31400 6812 -25480
rect 12732 -31400 12772 -25480
rect 6772 -31440 12772 -31400
rect 13384 -25480 19384 -25440
rect 13384 -31400 13424 -25480
rect 19344 -31400 19384 -25480
rect 13384 -31440 19384 -31400
rect 19996 -25480 25996 -25440
rect 19996 -31400 20036 -25480
rect 25956 -31400 25996 -25480
rect 19996 -31440 25996 -31400
rect 26608 -25480 32608 -25440
rect 26608 -31400 26648 -25480
rect 32568 -31400 32608 -25480
rect 26608 -31440 32608 -31400
rect 33220 -25480 39220 -25440
rect 33220 -31400 33260 -25480
rect 39180 -31400 39220 -25480
rect 33220 -31440 39220 -31400
rect -39512 -31800 -33512 -31760
rect -39512 -37720 -39472 -31800
rect -33552 -37720 -33512 -31800
rect -39512 -37760 -33512 -37720
rect -32900 -31800 -26900 -31760
rect -32900 -37720 -32860 -31800
rect -26940 -37720 -26900 -31800
rect -32900 -37760 -26900 -37720
rect -26288 -31800 -20288 -31760
rect -26288 -37720 -26248 -31800
rect -20328 -37720 -20288 -31800
rect -26288 -37760 -20288 -37720
rect -19676 -31800 -13676 -31760
rect -19676 -37720 -19636 -31800
rect -13716 -37720 -13676 -31800
rect -19676 -37760 -13676 -37720
rect -13064 -31800 -7064 -31760
rect -13064 -37720 -13024 -31800
rect -7104 -37720 -7064 -31800
rect -13064 -37760 -7064 -37720
rect -6452 -31800 -452 -31760
rect -6452 -37720 -6412 -31800
rect -492 -37720 -452 -31800
rect -6452 -37760 -452 -37720
rect 160 -31800 6160 -31760
rect 160 -37720 200 -31800
rect 6120 -37720 6160 -31800
rect 160 -37760 6160 -37720
rect 6772 -31800 12772 -31760
rect 6772 -37720 6812 -31800
rect 12732 -37720 12772 -31800
rect 6772 -37760 12772 -37720
rect 13384 -31800 19384 -31760
rect 13384 -37720 13424 -31800
rect 19344 -37720 19384 -31800
rect 13384 -37760 19384 -37720
rect 19996 -31800 25996 -31760
rect 19996 -37720 20036 -31800
rect 25956 -37720 25996 -31800
rect 19996 -37760 25996 -37720
rect 26608 -31800 32608 -31760
rect 26608 -37720 26648 -31800
rect 32568 -37720 32608 -31800
rect 26608 -37760 32608 -37720
rect 33220 -31800 39220 -31760
rect 33220 -37720 33260 -31800
rect 39180 -37720 39220 -31800
rect 33220 -37760 39220 -37720
<< mimcapcontact >>
rect -39472 31800 -33552 37720
rect -32860 31800 -26940 37720
rect -26248 31800 -20328 37720
rect -19636 31800 -13716 37720
rect -13024 31800 -7104 37720
rect -6412 31800 -492 37720
rect 200 31800 6120 37720
rect 6812 31800 12732 37720
rect 13424 31800 19344 37720
rect 20036 31800 25956 37720
rect 26648 31800 32568 37720
rect 33260 31800 39180 37720
rect -39472 25480 -33552 31400
rect -32860 25480 -26940 31400
rect -26248 25480 -20328 31400
rect -19636 25480 -13716 31400
rect -13024 25480 -7104 31400
rect -6412 25480 -492 31400
rect 200 25480 6120 31400
rect 6812 25480 12732 31400
rect 13424 25480 19344 31400
rect 20036 25480 25956 31400
rect 26648 25480 32568 31400
rect 33260 25480 39180 31400
rect -39472 19160 -33552 25080
rect -32860 19160 -26940 25080
rect -26248 19160 -20328 25080
rect -19636 19160 -13716 25080
rect -13024 19160 -7104 25080
rect -6412 19160 -492 25080
rect 200 19160 6120 25080
rect 6812 19160 12732 25080
rect 13424 19160 19344 25080
rect 20036 19160 25956 25080
rect 26648 19160 32568 25080
rect 33260 19160 39180 25080
rect -39472 12840 -33552 18760
rect -32860 12840 -26940 18760
rect -26248 12840 -20328 18760
rect -19636 12840 -13716 18760
rect -13024 12840 -7104 18760
rect -6412 12840 -492 18760
rect 200 12840 6120 18760
rect 6812 12840 12732 18760
rect 13424 12840 19344 18760
rect 20036 12840 25956 18760
rect 26648 12840 32568 18760
rect 33260 12840 39180 18760
rect -39472 6520 -33552 12440
rect -32860 6520 -26940 12440
rect -26248 6520 -20328 12440
rect -19636 6520 -13716 12440
rect -13024 6520 -7104 12440
rect -6412 6520 -492 12440
rect 200 6520 6120 12440
rect 6812 6520 12732 12440
rect 13424 6520 19344 12440
rect 20036 6520 25956 12440
rect 26648 6520 32568 12440
rect 33260 6520 39180 12440
rect -39472 200 -33552 6120
rect -32860 200 -26940 6120
rect -26248 200 -20328 6120
rect -19636 200 -13716 6120
rect -13024 200 -7104 6120
rect -6412 200 -492 6120
rect 200 200 6120 6120
rect 6812 200 12732 6120
rect 13424 200 19344 6120
rect 20036 200 25956 6120
rect 26648 200 32568 6120
rect 33260 200 39180 6120
rect -39472 -6120 -33552 -200
rect -32860 -6120 -26940 -200
rect -26248 -6120 -20328 -200
rect -19636 -6120 -13716 -200
rect -13024 -6120 -7104 -200
rect -6412 -6120 -492 -200
rect 200 -6120 6120 -200
rect 6812 -6120 12732 -200
rect 13424 -6120 19344 -200
rect 20036 -6120 25956 -200
rect 26648 -6120 32568 -200
rect 33260 -6120 39180 -200
rect -39472 -12440 -33552 -6520
rect -32860 -12440 -26940 -6520
rect -26248 -12440 -20328 -6520
rect -19636 -12440 -13716 -6520
rect -13024 -12440 -7104 -6520
rect -6412 -12440 -492 -6520
rect 200 -12440 6120 -6520
rect 6812 -12440 12732 -6520
rect 13424 -12440 19344 -6520
rect 20036 -12440 25956 -6520
rect 26648 -12440 32568 -6520
rect 33260 -12440 39180 -6520
rect -39472 -18760 -33552 -12840
rect -32860 -18760 -26940 -12840
rect -26248 -18760 -20328 -12840
rect -19636 -18760 -13716 -12840
rect -13024 -18760 -7104 -12840
rect -6412 -18760 -492 -12840
rect 200 -18760 6120 -12840
rect 6812 -18760 12732 -12840
rect 13424 -18760 19344 -12840
rect 20036 -18760 25956 -12840
rect 26648 -18760 32568 -12840
rect 33260 -18760 39180 -12840
rect -39472 -25080 -33552 -19160
rect -32860 -25080 -26940 -19160
rect -26248 -25080 -20328 -19160
rect -19636 -25080 -13716 -19160
rect -13024 -25080 -7104 -19160
rect -6412 -25080 -492 -19160
rect 200 -25080 6120 -19160
rect 6812 -25080 12732 -19160
rect 13424 -25080 19344 -19160
rect 20036 -25080 25956 -19160
rect 26648 -25080 32568 -19160
rect 33260 -25080 39180 -19160
rect -39472 -31400 -33552 -25480
rect -32860 -31400 -26940 -25480
rect -26248 -31400 -20328 -25480
rect -19636 -31400 -13716 -25480
rect -13024 -31400 -7104 -25480
rect -6412 -31400 -492 -25480
rect 200 -31400 6120 -25480
rect 6812 -31400 12732 -25480
rect 13424 -31400 19344 -25480
rect 20036 -31400 25956 -25480
rect 26648 -31400 32568 -25480
rect 33260 -31400 39180 -25480
rect -39472 -37720 -33552 -31800
rect -32860 -37720 -26940 -31800
rect -26248 -37720 -20328 -31800
rect -19636 -37720 -13716 -31800
rect -13024 -37720 -7104 -31800
rect -6412 -37720 -492 -31800
rect 200 -37720 6120 -31800
rect 6812 -37720 12732 -31800
rect 13424 -37720 19344 -31800
rect 20036 -37720 25956 -31800
rect 26648 -37720 32568 -31800
rect 33260 -37720 39180 -31800
<< metal4 >>
rect -36564 37721 -36460 37920
rect -33284 37772 -33180 37920
rect -39473 37720 -33551 37721
rect -39473 31800 -39472 37720
rect -33552 31800 -33551 37720
rect -39473 31799 -33551 31800
rect -36564 31401 -36460 31799
rect -33284 31748 -33264 37772
rect -33200 31748 -33180 37772
rect -29952 37721 -29848 37920
rect -26672 37772 -26568 37920
rect -32861 37720 -26939 37721
rect -32861 31800 -32860 37720
rect -26940 31800 -26939 37720
rect -32861 31799 -26939 31800
rect -33284 31452 -33180 31748
rect -39473 31400 -33551 31401
rect -39473 25480 -39472 31400
rect -33552 25480 -33551 31400
rect -39473 25479 -33551 25480
rect -36564 25081 -36460 25479
rect -33284 25428 -33264 31452
rect -33200 25428 -33180 31452
rect -29952 31401 -29848 31799
rect -26672 31748 -26652 37772
rect -26588 31748 -26568 37772
rect -23340 37721 -23236 37920
rect -20060 37772 -19956 37920
rect -26249 37720 -20327 37721
rect -26249 31800 -26248 37720
rect -20328 31800 -20327 37720
rect -26249 31799 -20327 31800
rect -26672 31452 -26568 31748
rect -32861 31400 -26939 31401
rect -32861 25480 -32860 31400
rect -26940 25480 -26939 31400
rect -32861 25479 -26939 25480
rect -33284 25132 -33180 25428
rect -39473 25080 -33551 25081
rect -39473 19160 -39472 25080
rect -33552 19160 -33551 25080
rect -39473 19159 -33551 19160
rect -36564 18761 -36460 19159
rect -33284 19108 -33264 25132
rect -33200 19108 -33180 25132
rect -29952 25081 -29848 25479
rect -26672 25428 -26652 31452
rect -26588 25428 -26568 31452
rect -23340 31401 -23236 31799
rect -20060 31748 -20040 37772
rect -19976 31748 -19956 37772
rect -16728 37721 -16624 37920
rect -13448 37772 -13344 37920
rect -19637 37720 -13715 37721
rect -19637 31800 -19636 37720
rect -13716 31800 -13715 37720
rect -19637 31799 -13715 31800
rect -20060 31452 -19956 31748
rect -26249 31400 -20327 31401
rect -26249 25480 -26248 31400
rect -20328 25480 -20327 31400
rect -26249 25479 -20327 25480
rect -26672 25132 -26568 25428
rect -32861 25080 -26939 25081
rect -32861 19160 -32860 25080
rect -26940 19160 -26939 25080
rect -32861 19159 -26939 19160
rect -33284 18812 -33180 19108
rect -39473 18760 -33551 18761
rect -39473 12840 -39472 18760
rect -33552 12840 -33551 18760
rect -39473 12839 -33551 12840
rect -36564 12441 -36460 12839
rect -33284 12788 -33264 18812
rect -33200 12788 -33180 18812
rect -29952 18761 -29848 19159
rect -26672 19108 -26652 25132
rect -26588 19108 -26568 25132
rect -23340 25081 -23236 25479
rect -20060 25428 -20040 31452
rect -19976 25428 -19956 31452
rect -16728 31401 -16624 31799
rect -13448 31748 -13428 37772
rect -13364 31748 -13344 37772
rect -10116 37721 -10012 37920
rect -6836 37772 -6732 37920
rect -13025 37720 -7103 37721
rect -13025 31800 -13024 37720
rect -7104 31800 -7103 37720
rect -13025 31799 -7103 31800
rect -13448 31452 -13344 31748
rect -19637 31400 -13715 31401
rect -19637 25480 -19636 31400
rect -13716 25480 -13715 31400
rect -19637 25479 -13715 25480
rect -20060 25132 -19956 25428
rect -26249 25080 -20327 25081
rect -26249 19160 -26248 25080
rect -20328 19160 -20327 25080
rect -26249 19159 -20327 19160
rect -26672 18812 -26568 19108
rect -32861 18760 -26939 18761
rect -32861 12840 -32860 18760
rect -26940 12840 -26939 18760
rect -32861 12839 -26939 12840
rect -33284 12492 -33180 12788
rect -39473 12440 -33551 12441
rect -39473 6520 -39472 12440
rect -33552 6520 -33551 12440
rect -39473 6519 -33551 6520
rect -36564 6121 -36460 6519
rect -33284 6468 -33264 12492
rect -33200 6468 -33180 12492
rect -29952 12441 -29848 12839
rect -26672 12788 -26652 18812
rect -26588 12788 -26568 18812
rect -23340 18761 -23236 19159
rect -20060 19108 -20040 25132
rect -19976 19108 -19956 25132
rect -16728 25081 -16624 25479
rect -13448 25428 -13428 31452
rect -13364 25428 -13344 31452
rect -10116 31401 -10012 31799
rect -6836 31748 -6816 37772
rect -6752 31748 -6732 37772
rect -3504 37721 -3400 37920
rect -224 37772 -120 37920
rect -6413 37720 -491 37721
rect -6413 31800 -6412 37720
rect -492 31800 -491 37720
rect -6413 31799 -491 31800
rect -6836 31452 -6732 31748
rect -13025 31400 -7103 31401
rect -13025 25480 -13024 31400
rect -7104 25480 -7103 31400
rect -13025 25479 -7103 25480
rect -13448 25132 -13344 25428
rect -19637 25080 -13715 25081
rect -19637 19160 -19636 25080
rect -13716 19160 -13715 25080
rect -19637 19159 -13715 19160
rect -20060 18812 -19956 19108
rect -26249 18760 -20327 18761
rect -26249 12840 -26248 18760
rect -20328 12840 -20327 18760
rect -26249 12839 -20327 12840
rect -26672 12492 -26568 12788
rect -32861 12440 -26939 12441
rect -32861 6520 -32860 12440
rect -26940 6520 -26939 12440
rect -32861 6519 -26939 6520
rect -33284 6172 -33180 6468
rect -39473 6120 -33551 6121
rect -39473 200 -39472 6120
rect -33552 200 -33551 6120
rect -39473 199 -33551 200
rect -36564 -199 -36460 199
rect -33284 148 -33264 6172
rect -33200 148 -33180 6172
rect -29952 6121 -29848 6519
rect -26672 6468 -26652 12492
rect -26588 6468 -26568 12492
rect -23340 12441 -23236 12839
rect -20060 12788 -20040 18812
rect -19976 12788 -19956 18812
rect -16728 18761 -16624 19159
rect -13448 19108 -13428 25132
rect -13364 19108 -13344 25132
rect -10116 25081 -10012 25479
rect -6836 25428 -6816 31452
rect -6752 25428 -6732 31452
rect -3504 31401 -3400 31799
rect -224 31748 -204 37772
rect -140 31748 -120 37772
rect 3108 37721 3212 37920
rect 6388 37772 6492 37920
rect 199 37720 6121 37721
rect 199 31800 200 37720
rect 6120 31800 6121 37720
rect 199 31799 6121 31800
rect -224 31452 -120 31748
rect -6413 31400 -491 31401
rect -6413 25480 -6412 31400
rect -492 25480 -491 31400
rect -6413 25479 -491 25480
rect -6836 25132 -6732 25428
rect -13025 25080 -7103 25081
rect -13025 19160 -13024 25080
rect -7104 19160 -7103 25080
rect -13025 19159 -7103 19160
rect -13448 18812 -13344 19108
rect -19637 18760 -13715 18761
rect -19637 12840 -19636 18760
rect -13716 12840 -13715 18760
rect -19637 12839 -13715 12840
rect -20060 12492 -19956 12788
rect -26249 12440 -20327 12441
rect -26249 6520 -26248 12440
rect -20328 6520 -20327 12440
rect -26249 6519 -20327 6520
rect -26672 6172 -26568 6468
rect -32861 6120 -26939 6121
rect -32861 200 -32860 6120
rect -26940 200 -26939 6120
rect -32861 199 -26939 200
rect -33284 -148 -33180 148
rect -39473 -200 -33551 -199
rect -39473 -6120 -39472 -200
rect -33552 -6120 -33551 -200
rect -39473 -6121 -33551 -6120
rect -36564 -6519 -36460 -6121
rect -33284 -6172 -33264 -148
rect -33200 -6172 -33180 -148
rect -29952 -199 -29848 199
rect -26672 148 -26652 6172
rect -26588 148 -26568 6172
rect -23340 6121 -23236 6519
rect -20060 6468 -20040 12492
rect -19976 6468 -19956 12492
rect -16728 12441 -16624 12839
rect -13448 12788 -13428 18812
rect -13364 12788 -13344 18812
rect -10116 18761 -10012 19159
rect -6836 19108 -6816 25132
rect -6752 19108 -6732 25132
rect -3504 25081 -3400 25479
rect -224 25428 -204 31452
rect -140 25428 -120 31452
rect 3108 31401 3212 31799
rect 6388 31748 6408 37772
rect 6472 31748 6492 37772
rect 9720 37721 9824 37920
rect 13000 37772 13104 37920
rect 6811 37720 12733 37721
rect 6811 31800 6812 37720
rect 12732 31800 12733 37720
rect 6811 31799 12733 31800
rect 6388 31452 6492 31748
rect 199 31400 6121 31401
rect 199 25480 200 31400
rect 6120 25480 6121 31400
rect 199 25479 6121 25480
rect -224 25132 -120 25428
rect -6413 25080 -491 25081
rect -6413 19160 -6412 25080
rect -492 19160 -491 25080
rect -6413 19159 -491 19160
rect -6836 18812 -6732 19108
rect -13025 18760 -7103 18761
rect -13025 12840 -13024 18760
rect -7104 12840 -7103 18760
rect -13025 12839 -7103 12840
rect -13448 12492 -13344 12788
rect -19637 12440 -13715 12441
rect -19637 6520 -19636 12440
rect -13716 6520 -13715 12440
rect -19637 6519 -13715 6520
rect -20060 6172 -19956 6468
rect -26249 6120 -20327 6121
rect -26249 200 -26248 6120
rect -20328 200 -20327 6120
rect -26249 199 -20327 200
rect -26672 -148 -26568 148
rect -32861 -200 -26939 -199
rect -32861 -6120 -32860 -200
rect -26940 -6120 -26939 -200
rect -32861 -6121 -26939 -6120
rect -33284 -6468 -33180 -6172
rect -39473 -6520 -33551 -6519
rect -39473 -12440 -39472 -6520
rect -33552 -12440 -33551 -6520
rect -39473 -12441 -33551 -12440
rect -36564 -12839 -36460 -12441
rect -33284 -12492 -33264 -6468
rect -33200 -12492 -33180 -6468
rect -29952 -6519 -29848 -6121
rect -26672 -6172 -26652 -148
rect -26588 -6172 -26568 -148
rect -23340 -199 -23236 199
rect -20060 148 -20040 6172
rect -19976 148 -19956 6172
rect -16728 6121 -16624 6519
rect -13448 6468 -13428 12492
rect -13364 6468 -13344 12492
rect -10116 12441 -10012 12839
rect -6836 12788 -6816 18812
rect -6752 12788 -6732 18812
rect -3504 18761 -3400 19159
rect -224 19108 -204 25132
rect -140 19108 -120 25132
rect 3108 25081 3212 25479
rect 6388 25428 6408 31452
rect 6472 25428 6492 31452
rect 9720 31401 9824 31799
rect 13000 31748 13020 37772
rect 13084 31748 13104 37772
rect 16332 37721 16436 37920
rect 19612 37772 19716 37920
rect 13423 37720 19345 37721
rect 13423 31800 13424 37720
rect 19344 31800 19345 37720
rect 13423 31799 19345 31800
rect 13000 31452 13104 31748
rect 6811 31400 12733 31401
rect 6811 25480 6812 31400
rect 12732 25480 12733 31400
rect 6811 25479 12733 25480
rect 6388 25132 6492 25428
rect 199 25080 6121 25081
rect 199 19160 200 25080
rect 6120 19160 6121 25080
rect 199 19159 6121 19160
rect -224 18812 -120 19108
rect -6413 18760 -491 18761
rect -6413 12840 -6412 18760
rect -492 12840 -491 18760
rect -6413 12839 -491 12840
rect -6836 12492 -6732 12788
rect -13025 12440 -7103 12441
rect -13025 6520 -13024 12440
rect -7104 6520 -7103 12440
rect -13025 6519 -7103 6520
rect -13448 6172 -13344 6468
rect -19637 6120 -13715 6121
rect -19637 200 -19636 6120
rect -13716 200 -13715 6120
rect -19637 199 -13715 200
rect -20060 -148 -19956 148
rect -26249 -200 -20327 -199
rect -26249 -6120 -26248 -200
rect -20328 -6120 -20327 -200
rect -26249 -6121 -20327 -6120
rect -26672 -6468 -26568 -6172
rect -32861 -6520 -26939 -6519
rect -32861 -12440 -32860 -6520
rect -26940 -12440 -26939 -6520
rect -32861 -12441 -26939 -12440
rect -33284 -12788 -33180 -12492
rect -39473 -12840 -33551 -12839
rect -39473 -18760 -39472 -12840
rect -33552 -18760 -33551 -12840
rect -39473 -18761 -33551 -18760
rect -36564 -19159 -36460 -18761
rect -33284 -18812 -33264 -12788
rect -33200 -18812 -33180 -12788
rect -29952 -12839 -29848 -12441
rect -26672 -12492 -26652 -6468
rect -26588 -12492 -26568 -6468
rect -23340 -6519 -23236 -6121
rect -20060 -6172 -20040 -148
rect -19976 -6172 -19956 -148
rect -16728 -199 -16624 199
rect -13448 148 -13428 6172
rect -13364 148 -13344 6172
rect -10116 6121 -10012 6519
rect -6836 6468 -6816 12492
rect -6752 6468 -6732 12492
rect -3504 12441 -3400 12839
rect -224 12788 -204 18812
rect -140 12788 -120 18812
rect 3108 18761 3212 19159
rect 6388 19108 6408 25132
rect 6472 19108 6492 25132
rect 9720 25081 9824 25479
rect 13000 25428 13020 31452
rect 13084 25428 13104 31452
rect 16332 31401 16436 31799
rect 19612 31748 19632 37772
rect 19696 31748 19716 37772
rect 22944 37721 23048 37920
rect 26224 37772 26328 37920
rect 20035 37720 25957 37721
rect 20035 31800 20036 37720
rect 25956 31800 25957 37720
rect 20035 31799 25957 31800
rect 19612 31452 19716 31748
rect 13423 31400 19345 31401
rect 13423 25480 13424 31400
rect 19344 25480 19345 31400
rect 13423 25479 19345 25480
rect 13000 25132 13104 25428
rect 6811 25080 12733 25081
rect 6811 19160 6812 25080
rect 12732 19160 12733 25080
rect 6811 19159 12733 19160
rect 6388 18812 6492 19108
rect 199 18760 6121 18761
rect 199 12840 200 18760
rect 6120 12840 6121 18760
rect 199 12839 6121 12840
rect -224 12492 -120 12788
rect -6413 12440 -491 12441
rect -6413 6520 -6412 12440
rect -492 6520 -491 12440
rect -6413 6519 -491 6520
rect -6836 6172 -6732 6468
rect -13025 6120 -7103 6121
rect -13025 200 -13024 6120
rect -7104 200 -7103 6120
rect -13025 199 -7103 200
rect -13448 -148 -13344 148
rect -19637 -200 -13715 -199
rect -19637 -6120 -19636 -200
rect -13716 -6120 -13715 -200
rect -19637 -6121 -13715 -6120
rect -20060 -6468 -19956 -6172
rect -26249 -6520 -20327 -6519
rect -26249 -12440 -26248 -6520
rect -20328 -12440 -20327 -6520
rect -26249 -12441 -20327 -12440
rect -26672 -12788 -26568 -12492
rect -32861 -12840 -26939 -12839
rect -32861 -18760 -32860 -12840
rect -26940 -18760 -26939 -12840
rect -32861 -18761 -26939 -18760
rect -33284 -19108 -33180 -18812
rect -39473 -19160 -33551 -19159
rect -39473 -25080 -39472 -19160
rect -33552 -25080 -33551 -19160
rect -39473 -25081 -33551 -25080
rect -36564 -25479 -36460 -25081
rect -33284 -25132 -33264 -19108
rect -33200 -25132 -33180 -19108
rect -29952 -19159 -29848 -18761
rect -26672 -18812 -26652 -12788
rect -26588 -18812 -26568 -12788
rect -23340 -12839 -23236 -12441
rect -20060 -12492 -20040 -6468
rect -19976 -12492 -19956 -6468
rect -16728 -6519 -16624 -6121
rect -13448 -6172 -13428 -148
rect -13364 -6172 -13344 -148
rect -10116 -199 -10012 199
rect -6836 148 -6816 6172
rect -6752 148 -6732 6172
rect -3504 6121 -3400 6519
rect -224 6468 -204 12492
rect -140 6468 -120 12492
rect 3108 12441 3212 12839
rect 6388 12788 6408 18812
rect 6472 12788 6492 18812
rect 9720 18761 9824 19159
rect 13000 19108 13020 25132
rect 13084 19108 13104 25132
rect 16332 25081 16436 25479
rect 19612 25428 19632 31452
rect 19696 25428 19716 31452
rect 22944 31401 23048 31799
rect 26224 31748 26244 37772
rect 26308 31748 26328 37772
rect 29556 37721 29660 37920
rect 32836 37772 32940 37920
rect 26647 37720 32569 37721
rect 26647 31800 26648 37720
rect 32568 31800 32569 37720
rect 26647 31799 32569 31800
rect 26224 31452 26328 31748
rect 20035 31400 25957 31401
rect 20035 25480 20036 31400
rect 25956 25480 25957 31400
rect 20035 25479 25957 25480
rect 19612 25132 19716 25428
rect 13423 25080 19345 25081
rect 13423 19160 13424 25080
rect 19344 19160 19345 25080
rect 13423 19159 19345 19160
rect 13000 18812 13104 19108
rect 6811 18760 12733 18761
rect 6811 12840 6812 18760
rect 12732 12840 12733 18760
rect 6811 12839 12733 12840
rect 6388 12492 6492 12788
rect 199 12440 6121 12441
rect 199 6520 200 12440
rect 6120 6520 6121 12440
rect 199 6519 6121 6520
rect -224 6172 -120 6468
rect -6413 6120 -491 6121
rect -6413 200 -6412 6120
rect -492 200 -491 6120
rect -6413 199 -491 200
rect -6836 -148 -6732 148
rect -13025 -200 -7103 -199
rect -13025 -6120 -13024 -200
rect -7104 -6120 -7103 -200
rect -13025 -6121 -7103 -6120
rect -13448 -6468 -13344 -6172
rect -19637 -6520 -13715 -6519
rect -19637 -12440 -19636 -6520
rect -13716 -12440 -13715 -6520
rect -19637 -12441 -13715 -12440
rect -20060 -12788 -19956 -12492
rect -26249 -12840 -20327 -12839
rect -26249 -18760 -26248 -12840
rect -20328 -18760 -20327 -12840
rect -26249 -18761 -20327 -18760
rect -26672 -19108 -26568 -18812
rect -32861 -19160 -26939 -19159
rect -32861 -25080 -32860 -19160
rect -26940 -25080 -26939 -19160
rect -32861 -25081 -26939 -25080
rect -33284 -25428 -33180 -25132
rect -39473 -25480 -33551 -25479
rect -39473 -31400 -39472 -25480
rect -33552 -31400 -33551 -25480
rect -39473 -31401 -33551 -31400
rect -36564 -31799 -36460 -31401
rect -33284 -31452 -33264 -25428
rect -33200 -31452 -33180 -25428
rect -29952 -25479 -29848 -25081
rect -26672 -25132 -26652 -19108
rect -26588 -25132 -26568 -19108
rect -23340 -19159 -23236 -18761
rect -20060 -18812 -20040 -12788
rect -19976 -18812 -19956 -12788
rect -16728 -12839 -16624 -12441
rect -13448 -12492 -13428 -6468
rect -13364 -12492 -13344 -6468
rect -10116 -6519 -10012 -6121
rect -6836 -6172 -6816 -148
rect -6752 -6172 -6732 -148
rect -3504 -199 -3400 199
rect -224 148 -204 6172
rect -140 148 -120 6172
rect 3108 6121 3212 6519
rect 6388 6468 6408 12492
rect 6472 6468 6492 12492
rect 9720 12441 9824 12839
rect 13000 12788 13020 18812
rect 13084 12788 13104 18812
rect 16332 18761 16436 19159
rect 19612 19108 19632 25132
rect 19696 19108 19716 25132
rect 22944 25081 23048 25479
rect 26224 25428 26244 31452
rect 26308 25428 26328 31452
rect 29556 31401 29660 31799
rect 32836 31748 32856 37772
rect 32920 31748 32940 37772
rect 36168 37721 36272 37920
rect 39448 37772 39552 37920
rect 33259 37720 39181 37721
rect 33259 31800 33260 37720
rect 39180 31800 39181 37720
rect 33259 31799 39181 31800
rect 32836 31452 32940 31748
rect 26647 31400 32569 31401
rect 26647 25480 26648 31400
rect 32568 25480 32569 31400
rect 26647 25479 32569 25480
rect 26224 25132 26328 25428
rect 20035 25080 25957 25081
rect 20035 19160 20036 25080
rect 25956 19160 25957 25080
rect 20035 19159 25957 19160
rect 19612 18812 19716 19108
rect 13423 18760 19345 18761
rect 13423 12840 13424 18760
rect 19344 12840 19345 18760
rect 13423 12839 19345 12840
rect 13000 12492 13104 12788
rect 6811 12440 12733 12441
rect 6811 6520 6812 12440
rect 12732 6520 12733 12440
rect 6811 6519 12733 6520
rect 6388 6172 6492 6468
rect 199 6120 6121 6121
rect 199 200 200 6120
rect 6120 200 6121 6120
rect 199 199 6121 200
rect -224 -148 -120 148
rect -6413 -200 -491 -199
rect -6413 -6120 -6412 -200
rect -492 -6120 -491 -200
rect -6413 -6121 -491 -6120
rect -6836 -6468 -6732 -6172
rect -13025 -6520 -7103 -6519
rect -13025 -12440 -13024 -6520
rect -7104 -12440 -7103 -6520
rect -13025 -12441 -7103 -12440
rect -13448 -12788 -13344 -12492
rect -19637 -12840 -13715 -12839
rect -19637 -18760 -19636 -12840
rect -13716 -18760 -13715 -12840
rect -19637 -18761 -13715 -18760
rect -20060 -19108 -19956 -18812
rect -26249 -19160 -20327 -19159
rect -26249 -25080 -26248 -19160
rect -20328 -25080 -20327 -19160
rect -26249 -25081 -20327 -25080
rect -26672 -25428 -26568 -25132
rect -32861 -25480 -26939 -25479
rect -32861 -31400 -32860 -25480
rect -26940 -31400 -26939 -25480
rect -32861 -31401 -26939 -31400
rect -33284 -31748 -33180 -31452
rect -39473 -31800 -33551 -31799
rect -39473 -37720 -39472 -31800
rect -33552 -37720 -33551 -31800
rect -39473 -37721 -33551 -37720
rect -36564 -37920 -36460 -37721
rect -33284 -37772 -33264 -31748
rect -33200 -37772 -33180 -31748
rect -29952 -31799 -29848 -31401
rect -26672 -31452 -26652 -25428
rect -26588 -31452 -26568 -25428
rect -23340 -25479 -23236 -25081
rect -20060 -25132 -20040 -19108
rect -19976 -25132 -19956 -19108
rect -16728 -19159 -16624 -18761
rect -13448 -18812 -13428 -12788
rect -13364 -18812 -13344 -12788
rect -10116 -12839 -10012 -12441
rect -6836 -12492 -6816 -6468
rect -6752 -12492 -6732 -6468
rect -3504 -6519 -3400 -6121
rect -224 -6172 -204 -148
rect -140 -6172 -120 -148
rect 3108 -199 3212 199
rect 6388 148 6408 6172
rect 6472 148 6492 6172
rect 9720 6121 9824 6519
rect 13000 6468 13020 12492
rect 13084 6468 13104 12492
rect 16332 12441 16436 12839
rect 19612 12788 19632 18812
rect 19696 12788 19716 18812
rect 22944 18761 23048 19159
rect 26224 19108 26244 25132
rect 26308 19108 26328 25132
rect 29556 25081 29660 25479
rect 32836 25428 32856 31452
rect 32920 25428 32940 31452
rect 36168 31401 36272 31799
rect 39448 31748 39468 37772
rect 39532 31748 39552 37772
rect 39448 31452 39552 31748
rect 33259 31400 39181 31401
rect 33259 25480 33260 31400
rect 39180 25480 39181 31400
rect 33259 25479 39181 25480
rect 32836 25132 32940 25428
rect 26647 25080 32569 25081
rect 26647 19160 26648 25080
rect 32568 19160 32569 25080
rect 26647 19159 32569 19160
rect 26224 18812 26328 19108
rect 20035 18760 25957 18761
rect 20035 12840 20036 18760
rect 25956 12840 25957 18760
rect 20035 12839 25957 12840
rect 19612 12492 19716 12788
rect 13423 12440 19345 12441
rect 13423 6520 13424 12440
rect 19344 6520 19345 12440
rect 13423 6519 19345 6520
rect 13000 6172 13104 6468
rect 6811 6120 12733 6121
rect 6811 200 6812 6120
rect 12732 200 12733 6120
rect 6811 199 12733 200
rect 6388 -148 6492 148
rect 199 -200 6121 -199
rect 199 -6120 200 -200
rect 6120 -6120 6121 -200
rect 199 -6121 6121 -6120
rect -224 -6468 -120 -6172
rect -6413 -6520 -491 -6519
rect -6413 -12440 -6412 -6520
rect -492 -12440 -491 -6520
rect -6413 -12441 -491 -12440
rect -6836 -12788 -6732 -12492
rect -13025 -12840 -7103 -12839
rect -13025 -18760 -13024 -12840
rect -7104 -18760 -7103 -12840
rect -13025 -18761 -7103 -18760
rect -13448 -19108 -13344 -18812
rect -19637 -19160 -13715 -19159
rect -19637 -25080 -19636 -19160
rect -13716 -25080 -13715 -19160
rect -19637 -25081 -13715 -25080
rect -20060 -25428 -19956 -25132
rect -26249 -25480 -20327 -25479
rect -26249 -31400 -26248 -25480
rect -20328 -31400 -20327 -25480
rect -26249 -31401 -20327 -31400
rect -26672 -31748 -26568 -31452
rect -32861 -31800 -26939 -31799
rect -32861 -37720 -32860 -31800
rect -26940 -37720 -26939 -31800
rect -32861 -37721 -26939 -37720
rect -33284 -37920 -33180 -37772
rect -29952 -37920 -29848 -37721
rect -26672 -37772 -26652 -31748
rect -26588 -37772 -26568 -31748
rect -23340 -31799 -23236 -31401
rect -20060 -31452 -20040 -25428
rect -19976 -31452 -19956 -25428
rect -16728 -25479 -16624 -25081
rect -13448 -25132 -13428 -19108
rect -13364 -25132 -13344 -19108
rect -10116 -19159 -10012 -18761
rect -6836 -18812 -6816 -12788
rect -6752 -18812 -6732 -12788
rect -3504 -12839 -3400 -12441
rect -224 -12492 -204 -6468
rect -140 -12492 -120 -6468
rect 3108 -6519 3212 -6121
rect 6388 -6172 6408 -148
rect 6472 -6172 6492 -148
rect 9720 -199 9824 199
rect 13000 148 13020 6172
rect 13084 148 13104 6172
rect 16332 6121 16436 6519
rect 19612 6468 19632 12492
rect 19696 6468 19716 12492
rect 22944 12441 23048 12839
rect 26224 12788 26244 18812
rect 26308 12788 26328 18812
rect 29556 18761 29660 19159
rect 32836 19108 32856 25132
rect 32920 19108 32940 25132
rect 36168 25081 36272 25479
rect 39448 25428 39468 31452
rect 39532 25428 39552 31452
rect 39448 25132 39552 25428
rect 33259 25080 39181 25081
rect 33259 19160 33260 25080
rect 39180 19160 39181 25080
rect 33259 19159 39181 19160
rect 32836 18812 32940 19108
rect 26647 18760 32569 18761
rect 26647 12840 26648 18760
rect 32568 12840 32569 18760
rect 26647 12839 32569 12840
rect 26224 12492 26328 12788
rect 20035 12440 25957 12441
rect 20035 6520 20036 12440
rect 25956 6520 25957 12440
rect 20035 6519 25957 6520
rect 19612 6172 19716 6468
rect 13423 6120 19345 6121
rect 13423 200 13424 6120
rect 19344 200 19345 6120
rect 13423 199 19345 200
rect 13000 -148 13104 148
rect 6811 -200 12733 -199
rect 6811 -6120 6812 -200
rect 12732 -6120 12733 -200
rect 6811 -6121 12733 -6120
rect 6388 -6468 6492 -6172
rect 199 -6520 6121 -6519
rect 199 -12440 200 -6520
rect 6120 -12440 6121 -6520
rect 199 -12441 6121 -12440
rect -224 -12788 -120 -12492
rect -6413 -12840 -491 -12839
rect -6413 -18760 -6412 -12840
rect -492 -18760 -491 -12840
rect -6413 -18761 -491 -18760
rect -6836 -19108 -6732 -18812
rect -13025 -19160 -7103 -19159
rect -13025 -25080 -13024 -19160
rect -7104 -25080 -7103 -19160
rect -13025 -25081 -7103 -25080
rect -13448 -25428 -13344 -25132
rect -19637 -25480 -13715 -25479
rect -19637 -31400 -19636 -25480
rect -13716 -31400 -13715 -25480
rect -19637 -31401 -13715 -31400
rect -20060 -31748 -19956 -31452
rect -26249 -31800 -20327 -31799
rect -26249 -37720 -26248 -31800
rect -20328 -37720 -20327 -31800
rect -26249 -37721 -20327 -37720
rect -26672 -37920 -26568 -37772
rect -23340 -37920 -23236 -37721
rect -20060 -37772 -20040 -31748
rect -19976 -37772 -19956 -31748
rect -16728 -31799 -16624 -31401
rect -13448 -31452 -13428 -25428
rect -13364 -31452 -13344 -25428
rect -10116 -25479 -10012 -25081
rect -6836 -25132 -6816 -19108
rect -6752 -25132 -6732 -19108
rect -3504 -19159 -3400 -18761
rect -224 -18812 -204 -12788
rect -140 -18812 -120 -12788
rect 3108 -12839 3212 -12441
rect 6388 -12492 6408 -6468
rect 6472 -12492 6492 -6468
rect 9720 -6519 9824 -6121
rect 13000 -6172 13020 -148
rect 13084 -6172 13104 -148
rect 16332 -199 16436 199
rect 19612 148 19632 6172
rect 19696 148 19716 6172
rect 22944 6121 23048 6519
rect 26224 6468 26244 12492
rect 26308 6468 26328 12492
rect 29556 12441 29660 12839
rect 32836 12788 32856 18812
rect 32920 12788 32940 18812
rect 36168 18761 36272 19159
rect 39448 19108 39468 25132
rect 39532 19108 39552 25132
rect 39448 18812 39552 19108
rect 33259 18760 39181 18761
rect 33259 12840 33260 18760
rect 39180 12840 39181 18760
rect 33259 12839 39181 12840
rect 32836 12492 32940 12788
rect 26647 12440 32569 12441
rect 26647 6520 26648 12440
rect 32568 6520 32569 12440
rect 26647 6519 32569 6520
rect 26224 6172 26328 6468
rect 20035 6120 25957 6121
rect 20035 200 20036 6120
rect 25956 200 25957 6120
rect 20035 199 25957 200
rect 19612 -148 19716 148
rect 13423 -200 19345 -199
rect 13423 -6120 13424 -200
rect 19344 -6120 19345 -200
rect 13423 -6121 19345 -6120
rect 13000 -6468 13104 -6172
rect 6811 -6520 12733 -6519
rect 6811 -12440 6812 -6520
rect 12732 -12440 12733 -6520
rect 6811 -12441 12733 -12440
rect 6388 -12788 6492 -12492
rect 199 -12840 6121 -12839
rect 199 -18760 200 -12840
rect 6120 -18760 6121 -12840
rect 199 -18761 6121 -18760
rect -224 -19108 -120 -18812
rect -6413 -19160 -491 -19159
rect -6413 -25080 -6412 -19160
rect -492 -25080 -491 -19160
rect -6413 -25081 -491 -25080
rect -6836 -25428 -6732 -25132
rect -13025 -25480 -7103 -25479
rect -13025 -31400 -13024 -25480
rect -7104 -31400 -7103 -25480
rect -13025 -31401 -7103 -31400
rect -13448 -31748 -13344 -31452
rect -19637 -31800 -13715 -31799
rect -19637 -37720 -19636 -31800
rect -13716 -37720 -13715 -31800
rect -19637 -37721 -13715 -37720
rect -20060 -37920 -19956 -37772
rect -16728 -37920 -16624 -37721
rect -13448 -37772 -13428 -31748
rect -13364 -37772 -13344 -31748
rect -10116 -31799 -10012 -31401
rect -6836 -31452 -6816 -25428
rect -6752 -31452 -6732 -25428
rect -3504 -25479 -3400 -25081
rect -224 -25132 -204 -19108
rect -140 -25132 -120 -19108
rect 3108 -19159 3212 -18761
rect 6388 -18812 6408 -12788
rect 6472 -18812 6492 -12788
rect 9720 -12839 9824 -12441
rect 13000 -12492 13020 -6468
rect 13084 -12492 13104 -6468
rect 16332 -6519 16436 -6121
rect 19612 -6172 19632 -148
rect 19696 -6172 19716 -148
rect 22944 -199 23048 199
rect 26224 148 26244 6172
rect 26308 148 26328 6172
rect 29556 6121 29660 6519
rect 32836 6468 32856 12492
rect 32920 6468 32940 12492
rect 36168 12441 36272 12839
rect 39448 12788 39468 18812
rect 39532 12788 39552 18812
rect 39448 12492 39552 12788
rect 33259 12440 39181 12441
rect 33259 6520 33260 12440
rect 39180 6520 39181 12440
rect 33259 6519 39181 6520
rect 32836 6172 32940 6468
rect 26647 6120 32569 6121
rect 26647 200 26648 6120
rect 32568 200 32569 6120
rect 26647 199 32569 200
rect 26224 -148 26328 148
rect 20035 -200 25957 -199
rect 20035 -6120 20036 -200
rect 25956 -6120 25957 -200
rect 20035 -6121 25957 -6120
rect 19612 -6468 19716 -6172
rect 13423 -6520 19345 -6519
rect 13423 -12440 13424 -6520
rect 19344 -12440 19345 -6520
rect 13423 -12441 19345 -12440
rect 13000 -12788 13104 -12492
rect 6811 -12840 12733 -12839
rect 6811 -18760 6812 -12840
rect 12732 -18760 12733 -12840
rect 6811 -18761 12733 -18760
rect 6388 -19108 6492 -18812
rect 199 -19160 6121 -19159
rect 199 -25080 200 -19160
rect 6120 -25080 6121 -19160
rect 199 -25081 6121 -25080
rect -224 -25428 -120 -25132
rect -6413 -25480 -491 -25479
rect -6413 -31400 -6412 -25480
rect -492 -31400 -491 -25480
rect -6413 -31401 -491 -31400
rect -6836 -31748 -6732 -31452
rect -13025 -31800 -7103 -31799
rect -13025 -37720 -13024 -31800
rect -7104 -37720 -7103 -31800
rect -13025 -37721 -7103 -37720
rect -13448 -37920 -13344 -37772
rect -10116 -37920 -10012 -37721
rect -6836 -37772 -6816 -31748
rect -6752 -37772 -6732 -31748
rect -3504 -31799 -3400 -31401
rect -224 -31452 -204 -25428
rect -140 -31452 -120 -25428
rect 3108 -25479 3212 -25081
rect 6388 -25132 6408 -19108
rect 6472 -25132 6492 -19108
rect 9720 -19159 9824 -18761
rect 13000 -18812 13020 -12788
rect 13084 -18812 13104 -12788
rect 16332 -12839 16436 -12441
rect 19612 -12492 19632 -6468
rect 19696 -12492 19716 -6468
rect 22944 -6519 23048 -6121
rect 26224 -6172 26244 -148
rect 26308 -6172 26328 -148
rect 29556 -199 29660 199
rect 32836 148 32856 6172
rect 32920 148 32940 6172
rect 36168 6121 36272 6519
rect 39448 6468 39468 12492
rect 39532 6468 39552 12492
rect 39448 6172 39552 6468
rect 33259 6120 39181 6121
rect 33259 200 33260 6120
rect 39180 200 39181 6120
rect 33259 199 39181 200
rect 32836 -148 32940 148
rect 26647 -200 32569 -199
rect 26647 -6120 26648 -200
rect 32568 -6120 32569 -200
rect 26647 -6121 32569 -6120
rect 26224 -6468 26328 -6172
rect 20035 -6520 25957 -6519
rect 20035 -12440 20036 -6520
rect 25956 -12440 25957 -6520
rect 20035 -12441 25957 -12440
rect 19612 -12788 19716 -12492
rect 13423 -12840 19345 -12839
rect 13423 -18760 13424 -12840
rect 19344 -18760 19345 -12840
rect 13423 -18761 19345 -18760
rect 13000 -19108 13104 -18812
rect 6811 -19160 12733 -19159
rect 6811 -25080 6812 -19160
rect 12732 -25080 12733 -19160
rect 6811 -25081 12733 -25080
rect 6388 -25428 6492 -25132
rect 199 -25480 6121 -25479
rect 199 -31400 200 -25480
rect 6120 -31400 6121 -25480
rect 199 -31401 6121 -31400
rect -224 -31748 -120 -31452
rect -6413 -31800 -491 -31799
rect -6413 -37720 -6412 -31800
rect -492 -37720 -491 -31800
rect -6413 -37721 -491 -37720
rect -6836 -37920 -6732 -37772
rect -3504 -37920 -3400 -37721
rect -224 -37772 -204 -31748
rect -140 -37772 -120 -31748
rect 3108 -31799 3212 -31401
rect 6388 -31452 6408 -25428
rect 6472 -31452 6492 -25428
rect 9720 -25479 9824 -25081
rect 13000 -25132 13020 -19108
rect 13084 -25132 13104 -19108
rect 16332 -19159 16436 -18761
rect 19612 -18812 19632 -12788
rect 19696 -18812 19716 -12788
rect 22944 -12839 23048 -12441
rect 26224 -12492 26244 -6468
rect 26308 -12492 26328 -6468
rect 29556 -6519 29660 -6121
rect 32836 -6172 32856 -148
rect 32920 -6172 32940 -148
rect 36168 -199 36272 199
rect 39448 148 39468 6172
rect 39532 148 39552 6172
rect 39448 -148 39552 148
rect 33259 -200 39181 -199
rect 33259 -6120 33260 -200
rect 39180 -6120 39181 -200
rect 33259 -6121 39181 -6120
rect 32836 -6468 32940 -6172
rect 26647 -6520 32569 -6519
rect 26647 -12440 26648 -6520
rect 32568 -12440 32569 -6520
rect 26647 -12441 32569 -12440
rect 26224 -12788 26328 -12492
rect 20035 -12840 25957 -12839
rect 20035 -18760 20036 -12840
rect 25956 -18760 25957 -12840
rect 20035 -18761 25957 -18760
rect 19612 -19108 19716 -18812
rect 13423 -19160 19345 -19159
rect 13423 -25080 13424 -19160
rect 19344 -25080 19345 -19160
rect 13423 -25081 19345 -25080
rect 13000 -25428 13104 -25132
rect 6811 -25480 12733 -25479
rect 6811 -31400 6812 -25480
rect 12732 -31400 12733 -25480
rect 6811 -31401 12733 -31400
rect 6388 -31748 6492 -31452
rect 199 -31800 6121 -31799
rect 199 -37720 200 -31800
rect 6120 -37720 6121 -31800
rect 199 -37721 6121 -37720
rect -224 -37920 -120 -37772
rect 3108 -37920 3212 -37721
rect 6388 -37772 6408 -31748
rect 6472 -37772 6492 -31748
rect 9720 -31799 9824 -31401
rect 13000 -31452 13020 -25428
rect 13084 -31452 13104 -25428
rect 16332 -25479 16436 -25081
rect 19612 -25132 19632 -19108
rect 19696 -25132 19716 -19108
rect 22944 -19159 23048 -18761
rect 26224 -18812 26244 -12788
rect 26308 -18812 26328 -12788
rect 29556 -12839 29660 -12441
rect 32836 -12492 32856 -6468
rect 32920 -12492 32940 -6468
rect 36168 -6519 36272 -6121
rect 39448 -6172 39468 -148
rect 39532 -6172 39552 -148
rect 39448 -6468 39552 -6172
rect 33259 -6520 39181 -6519
rect 33259 -12440 33260 -6520
rect 39180 -12440 39181 -6520
rect 33259 -12441 39181 -12440
rect 32836 -12788 32940 -12492
rect 26647 -12840 32569 -12839
rect 26647 -18760 26648 -12840
rect 32568 -18760 32569 -12840
rect 26647 -18761 32569 -18760
rect 26224 -19108 26328 -18812
rect 20035 -19160 25957 -19159
rect 20035 -25080 20036 -19160
rect 25956 -25080 25957 -19160
rect 20035 -25081 25957 -25080
rect 19612 -25428 19716 -25132
rect 13423 -25480 19345 -25479
rect 13423 -31400 13424 -25480
rect 19344 -31400 19345 -25480
rect 13423 -31401 19345 -31400
rect 13000 -31748 13104 -31452
rect 6811 -31800 12733 -31799
rect 6811 -37720 6812 -31800
rect 12732 -37720 12733 -31800
rect 6811 -37721 12733 -37720
rect 6388 -37920 6492 -37772
rect 9720 -37920 9824 -37721
rect 13000 -37772 13020 -31748
rect 13084 -37772 13104 -31748
rect 16332 -31799 16436 -31401
rect 19612 -31452 19632 -25428
rect 19696 -31452 19716 -25428
rect 22944 -25479 23048 -25081
rect 26224 -25132 26244 -19108
rect 26308 -25132 26328 -19108
rect 29556 -19159 29660 -18761
rect 32836 -18812 32856 -12788
rect 32920 -18812 32940 -12788
rect 36168 -12839 36272 -12441
rect 39448 -12492 39468 -6468
rect 39532 -12492 39552 -6468
rect 39448 -12788 39552 -12492
rect 33259 -12840 39181 -12839
rect 33259 -18760 33260 -12840
rect 39180 -18760 39181 -12840
rect 33259 -18761 39181 -18760
rect 32836 -19108 32940 -18812
rect 26647 -19160 32569 -19159
rect 26647 -25080 26648 -19160
rect 32568 -25080 32569 -19160
rect 26647 -25081 32569 -25080
rect 26224 -25428 26328 -25132
rect 20035 -25480 25957 -25479
rect 20035 -31400 20036 -25480
rect 25956 -31400 25957 -25480
rect 20035 -31401 25957 -31400
rect 19612 -31748 19716 -31452
rect 13423 -31800 19345 -31799
rect 13423 -37720 13424 -31800
rect 19344 -37720 19345 -31800
rect 13423 -37721 19345 -37720
rect 13000 -37920 13104 -37772
rect 16332 -37920 16436 -37721
rect 19612 -37772 19632 -31748
rect 19696 -37772 19716 -31748
rect 22944 -31799 23048 -31401
rect 26224 -31452 26244 -25428
rect 26308 -31452 26328 -25428
rect 29556 -25479 29660 -25081
rect 32836 -25132 32856 -19108
rect 32920 -25132 32940 -19108
rect 36168 -19159 36272 -18761
rect 39448 -18812 39468 -12788
rect 39532 -18812 39552 -12788
rect 39448 -19108 39552 -18812
rect 33259 -19160 39181 -19159
rect 33259 -25080 33260 -19160
rect 39180 -25080 39181 -19160
rect 33259 -25081 39181 -25080
rect 32836 -25428 32940 -25132
rect 26647 -25480 32569 -25479
rect 26647 -31400 26648 -25480
rect 32568 -31400 32569 -25480
rect 26647 -31401 32569 -31400
rect 26224 -31748 26328 -31452
rect 20035 -31800 25957 -31799
rect 20035 -37720 20036 -31800
rect 25956 -37720 25957 -31800
rect 20035 -37721 25957 -37720
rect 19612 -37920 19716 -37772
rect 22944 -37920 23048 -37721
rect 26224 -37772 26244 -31748
rect 26308 -37772 26328 -31748
rect 29556 -31799 29660 -31401
rect 32836 -31452 32856 -25428
rect 32920 -31452 32940 -25428
rect 36168 -25479 36272 -25081
rect 39448 -25132 39468 -19108
rect 39532 -25132 39552 -19108
rect 39448 -25428 39552 -25132
rect 33259 -25480 39181 -25479
rect 33259 -31400 33260 -25480
rect 39180 -31400 39181 -25480
rect 33259 -31401 39181 -31400
rect 32836 -31748 32940 -31452
rect 26647 -31800 32569 -31799
rect 26647 -37720 26648 -31800
rect 32568 -37720 32569 -31800
rect 26647 -37721 32569 -37720
rect 26224 -37920 26328 -37772
rect 29556 -37920 29660 -37721
rect 32836 -37772 32856 -31748
rect 32920 -37772 32940 -31748
rect 36168 -31799 36272 -31401
rect 39448 -31452 39468 -25428
rect 39532 -31452 39552 -25428
rect 39448 -31748 39552 -31452
rect 33259 -31800 39181 -31799
rect 33259 -37720 33260 -31800
rect 39180 -37720 39181 -31800
rect 33259 -37721 39181 -37720
rect 32836 -37920 32940 -37772
rect 36168 -37920 36272 -37721
rect 39448 -37772 39468 -31748
rect 39532 -37772 39552 -31748
rect 39448 -37920 39552 -37772
<< properties >>
string FIXED_BBOX 33180 31720 39260 37800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 12 ny 12 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
