magic
tech sky130A
magscale 1 2
timestamp 1714283992
<< pwell >>
rect -214 -761 214 761
<< psubdiff >>
rect -178 691 -82 725
rect 82 691 178 725
rect -178 629 -144 691
rect 144 629 178 691
rect -178 -691 -144 -629
rect 144 -691 178 -629
rect -178 -725 -82 -691
rect 82 -725 178 -691
<< psubdiffcont >>
rect -82 691 82 725
rect -178 -629 -144 629
rect 144 -629 178 629
rect -82 -725 82 -691
<< poly >>
rect -48 579 48 595
rect -48 545 -32 579
rect 32 545 48 579
rect -48 165 48 545
rect -48 -545 48 -165
rect -48 -579 -32 -545
rect 32 -579 48 -545
rect -48 -595 48 -579
<< polycont >>
rect -32 545 32 579
rect -32 -579 32 -545
<< npolyres >>
rect -48 -165 48 165
<< locali >>
rect -178 691 -82 725
rect 82 691 178 725
rect -178 629 -144 691
rect 144 629 178 691
rect -48 545 -32 579
rect 32 545 48 579
rect -48 -579 -32 -545
rect 32 -579 48 -545
rect -178 -691 -144 -629
rect 144 -691 178 -629
rect -178 -725 -82 -691
rect 82 -725 178 -691
<< viali >>
rect -32 545 32 579
rect -32 182 32 545
rect -32 -545 32 -182
rect -32 -579 32 -545
<< metal1 >>
rect -38 579 38 591
rect -38 182 -32 579
rect 32 182 38 579
rect -38 170 38 182
rect -38 -182 38 -170
rect -38 -579 -32 -182
rect 32 -579 38 -182
rect -38 -591 38 -579
<< properties >>
string FIXED_BBOX -161 -708 161 708
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.48 l 1.650 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 165.687 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
