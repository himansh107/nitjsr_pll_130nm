magic
tech sky130A
magscale 1 2
timestamp 1714832304
<< metal1 >>
rect 17418 5002 18360 5070
rect 8859 3799 11051 3865
rect 11117 3799 11123 3865
rect 16801 3673 17211 3731
rect 11045 3275 11051 3341
rect 11117 3275 11123 3341
rect 11051 3200 11117 3275
rect -1669 3081 -58 3151
rect -1669 2605 -1599 3081
rect 11038 2952 12314 3200
rect 11051 2725 11117 2952
rect 11051 2653 11117 2659
rect 16240 2358 16560 2446
rect 16648 2358 16654 2446
rect -6340 2146 -6018 2196
rect 9710 1224 9778 1842
rect 8878 1156 8884 1224
rect 8952 1156 9778 1224
rect 10281 1785 11051 1851
rect 11117 1785 11123 1851
rect 8878 698 8884 766
rect 8952 698 8958 766
rect -6235 -2107 -6169 -461
rect -1567 -767 295 -705
rect 8884 -1756 8952 698
rect 10281 -19 10347 1785
rect 16801 589 16859 3673
rect 17426 852 17494 5002
rect 17690 2446 17778 2452
rect 17778 2358 18326 2446
rect 17690 2352 17778 2358
rect 17426 784 21494 852
rect 16801 531 20595 589
rect 20537 295 20595 531
rect 21426 416 21494 784
rect 22876 822 23204 888
rect 21426 342 21494 348
rect 22512 295 22628 674
rect 20537 237 22628 295
rect 21420 114 21426 182
rect 21494 114 21500 182
rect 21426 12 21494 114
rect 22570 -1066 22628 237
rect -6235 -2173 1141 -2107
rect 9616 -2120 9684 -2114
rect 1075 -3581 1141 -2173
rect 8200 -2188 9294 -2120
rect 9362 -2188 9368 -2120
rect 9684 -2188 9878 -2120
rect 9616 -2194 9684 -2188
rect 8202 -3062 8788 -2858
rect 22876 -3581 22942 822
rect 1075 -3647 22942 -3581
<< via1 >>
rect 11051 3799 11117 3865
rect 11051 3275 11117 3341
rect 11051 2659 11117 2725
rect 16560 2358 16648 2446
rect 8884 1156 8952 1224
rect 11051 1785 11117 1851
rect 8884 698 8952 766
rect 17690 2358 17778 2446
rect 21426 348 21494 416
rect 21426 114 21494 182
rect 9294 -2188 9362 -2120
rect 9616 -2188 9684 -2120
<< metal2 >>
rect 11051 3865 11117 3871
rect 11051 3341 11117 3799
rect 11051 3269 11117 3275
rect 11045 2659 11051 2725
rect 11117 2659 11123 2725
rect 11051 1851 11117 2659
rect 16560 2446 16648 2452
rect 16648 2358 17690 2446
rect 17778 2358 17784 2446
rect 16560 2352 16648 2358
rect 11051 1779 11117 1785
rect 8884 1224 8952 1230
rect 8884 766 8952 1156
rect 8884 692 8952 698
rect 21420 348 21426 416
rect 21494 348 21500 416
rect 21426 182 21494 348
rect 21426 108 21494 114
rect 9294 -2120 9362 -2114
rect 9362 -2188 9616 -2120
rect 9684 -2188 9690 -2120
rect 9294 -2194 9362 -2188
use cp  cp_0
timestamp 1714832304
transform 1 0 622 0 1 -2316
box -65526 -1044 51767 88502
use pfd_lay  pfd_lay_0
timestamp 1714832304
transform 1 0 -6940 0 1 1602
box 650 -3176 7450 1322
<< labels >>
flabel metal1 12148 3064 12148 3064 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel metal1 8664 -2964 8664 -2964 0 FreeSans 1600 0 0 0 GND
port 3 nsew
flabel metal1 -6312 2170 -6312 2170 0 FreeSans 480 0 0 0 f_clk_in
port 5 nsew
flabel metal1 22554 596 22554 596 0 FreeSans 480 0 0 0 f_clk_out
port 7 nsew
<< end >>
